(* blackbox *)
module qubitbytes_logo (
`ifdef USE_POWER_PINS
    input  VPWR,
    input  VGND
`endif  // USE_POWER_PINS
);
endmodule
