(* blackbox *)
module qubitbytes_logo (
`ifdef USE_POWER_PINS
    input  VGND,
    input  VPWR
`endif  // USE_POWER_PINS
);
endmodule
