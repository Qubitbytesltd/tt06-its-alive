VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO qubitbytes_logo
  CLASS BLOCK ;
  FOREIGN qubitbytes_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END qubitbytes_logo
END LIBRARY

