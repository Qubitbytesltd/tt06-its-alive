VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO qubitbytes_logo
  CLASS BLOCK ;
  FOREIGN qubitbytes_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.000 24.000 1.500 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 54.500 0.000 78.500 1.500 ;
    END
  END VGND
  OBS
      LAYER met1 ;
        RECT 0.000 9.500 78.500 25.500 ;
      LAYER met2 ;
        RECT 0.000 9.500 78.500 25.500 ;
      LAYER met3 ;
        RECT 0.000 9.500 78.500 25.500 ;
      LAYER met4 ;
        RECT 0.000 24.100 78.500 25.500 ;
        RECT 0.000 23.300 5.200 24.100 ;
      LAYER met4 ;
        RECT 5.200 23.300 11.600 24.100 ;
      LAYER met4 ;
        RECT 11.600 23.300 15.600 24.100 ;
      LAYER met4 ;
        RECT 15.600 23.300 16.400 24.100 ;
      LAYER met4 ;
        RECT 16.400 23.300 19.600 24.100 ;
      LAYER met4 ;
        RECT 19.600 23.300 20.400 24.100 ;
      LAYER met4 ;
        RECT 20.400 23.300 22.000 24.100 ;
        RECT 0.000 22.500 4.400 23.300 ;
      LAYER met4 ;
        RECT 4.400 22.500 11.600 23.300 ;
      LAYER met4 ;
        RECT 11.600 22.500 14.800 23.300 ;
      LAYER met4 ;
        RECT 14.800 22.500 16.400 23.300 ;
      LAYER met4 ;
        RECT 16.400 22.500 18.800 23.300 ;
      LAYER met4 ;
        RECT 18.800 22.500 21.200 23.300 ;
      LAYER met4 ;
        RECT 0.000 17.700 3.600 22.500 ;
      LAYER met4 ;
        RECT 3.600 17.700 6.000 22.500 ;
      LAYER met4 ;
        RECT 6.000 19.300 9.200 22.500 ;
      LAYER met4 ;
        RECT 9.200 20.900 11.600 22.500 ;
      LAYER met4 ;
        RECT 11.600 20.900 14.000 22.500 ;
      LAYER met4 ;
        RECT 9.200 20.100 10.800 20.900 ;
      LAYER met4 ;
        RECT 10.800 20.100 14.000 20.900 ;
      LAYER met4 ;
        RECT 9.200 19.300 10.000 20.100 ;
      LAYER met4 ;
        RECT 10.000 19.300 14.000 20.100 ;
      LAYER met4 ;
        RECT 14.000 19.300 16.400 22.500 ;
      LAYER met4 ;
        RECT 16.400 21.700 18.000 22.500 ;
      LAYER met4 ;
        RECT 18.000 21.700 21.200 22.500 ;
      LAYER met4 ;
        RECT 21.200 21.700 22.000 23.300 ;
        RECT 16.400 19.300 17.200 21.700 ;
      LAYER met4 ;
        RECT 17.200 20.900 20.400 21.700 ;
      LAYER met4 ;
        RECT 20.400 20.900 22.000 21.700 ;
      LAYER met4 ;
        RECT 17.200 20.100 19.600 20.900 ;
      LAYER met4 ;
        RECT 19.600 20.100 22.000 20.900 ;
      LAYER met4 ;
        RECT 17.200 19.300 18.800 20.100 ;
      LAYER met4 ;
        RECT 6.000 18.500 14.000 19.300 ;
      LAYER met4 ;
        RECT 14.000 18.500 18.800 19.300 ;
      LAYER met4 ;
        RECT 18.800 18.500 22.000 20.100 ;
        RECT 6.000 17.700 13.200 18.500 ;
      LAYER met4 ;
        RECT 13.200 17.700 18.000 18.500 ;
      LAYER met4 ;
        RECT 0.000 16.900 2.000 17.700 ;
      LAYER met4 ;
        RECT 2.000 16.900 11.600 17.700 ;
      LAYER met4 ;
        RECT 11.600 16.900 12.400 17.700 ;
      LAYER met4 ;
        RECT 12.400 16.900 18.000 17.700 ;
      LAYER met4 ;
        RECT 18.000 16.900 22.000 18.500 ;
        RECT 0.000 16.100 2.800 16.900 ;
      LAYER met4 ;
        RECT 2.800 16.100 11.600 16.900 ;
      LAYER met4 ;
        RECT 0.000 14.500 9.200 16.100 ;
        RECT 0.000 13.700 5.200 14.500 ;
      LAYER met4 ;
        RECT 5.200 13.700 6.000 14.500 ;
      LAYER met4 ;
        RECT 0.000 12.900 4.400 13.700 ;
      LAYER met4 ;
        RECT 4.400 12.900 6.000 13.700 ;
      LAYER met4 ;
        RECT 6.000 12.900 9.200 14.500 ;
      LAYER met4 ;
        RECT 9.200 12.900 11.600 16.100 ;
      LAYER met4 ;
        RECT 11.600 12.900 14.000 16.900 ;
      LAYER met4 ;
        RECT 14.000 16.100 18.800 16.900 ;
      LAYER met4 ;
        RECT 0.000 12.100 3.600 12.900 ;
      LAYER met4 ;
        RECT 3.600 12.100 10.800 12.900 ;
      LAYER met4 ;
        RECT 10.800 12.100 14.000 12.900 ;
        RECT 0.000 11.300 2.800 12.100 ;
      LAYER met4 ;
        RECT 2.800 11.300 10.000 12.100 ;
      LAYER met4 ;
        RECT 10.000 11.300 14.000 12.100 ;
      LAYER met4 ;
        RECT 14.000 11.300 16.400 16.100 ;
      LAYER met4 ;
        RECT 16.400 13.700 17.200 16.100 ;
      LAYER met4 ;
        RECT 17.200 15.300 18.800 16.100 ;
      LAYER met4 ;
        RECT 18.800 15.300 22.000 16.900 ;
      LAYER met4 ;
        RECT 17.200 14.500 19.600 15.300 ;
      LAYER met4 ;
        RECT 19.600 14.500 22.000 15.300 ;
      LAYER met4 ;
        RECT 17.200 13.700 20.400 14.500 ;
      LAYER met4 ;
        RECT 20.400 13.700 22.000 14.500 ;
        RECT 16.400 12.900 18.000 13.700 ;
      LAYER met4 ;
        RECT 18.000 12.900 21.200 13.700 ;
      LAYER met4 ;
        RECT 16.400 12.100 18.800 12.900 ;
      LAYER met4 ;
        RECT 18.800 12.100 21.200 12.900 ;
      LAYER met4 ;
        RECT 21.200 12.100 22.000 13.700 ;
      LAYER met4 ;
        RECT 22.000 12.900 24.400 24.100 ;
      LAYER met4 ;
        RECT 24.400 12.900 27.600 24.100 ;
      LAYER met4 ;
        RECT 27.600 23.300 28.400 24.100 ;
      LAYER met4 ;
        RECT 28.400 23.300 32.400 24.100 ;
      LAYER met4 ;
        RECT 32.400 23.300 33.200 24.100 ;
      LAYER met4 ;
        RECT 33.200 23.300 40.400 24.100 ;
      LAYER met4 ;
        RECT 40.400 23.300 41.200 24.100 ;
      LAYER met4 ;
        RECT 41.200 23.300 50.000 24.100 ;
      LAYER met4 ;
        RECT 50.000 23.300 56.400 24.100 ;
      LAYER met4 ;
        RECT 56.400 23.300 60.400 24.100 ;
      LAYER met4 ;
        RECT 60.400 23.300 66.800 24.100 ;
        RECT 27.600 22.500 29.200 23.300 ;
      LAYER met4 ;
        RECT 29.200 22.500 31.600 23.300 ;
      LAYER met4 ;
        RECT 31.600 22.500 33.200 23.300 ;
      LAYER met4 ;
        RECT 33.200 22.500 39.600 23.300 ;
      LAYER met4 ;
        RECT 39.600 22.500 41.200 23.300 ;
      LAYER met4 ;
        RECT 41.200 22.500 49.200 23.300 ;
      LAYER met4 ;
        RECT 49.200 22.500 56.400 23.300 ;
      LAYER met4 ;
        RECT 56.400 22.500 59.600 23.300 ;
      LAYER met4 ;
        RECT 59.600 22.500 66.800 23.300 ;
      LAYER met4 ;
        RECT 66.800 22.500 70.800 24.100 ;
      LAYER met4 ;
        RECT 70.800 22.500 73.200 24.100 ;
      LAYER met4 ;
        RECT 73.200 22.500 78.500 24.100 ;
      LAYER met4 ;
        RECT 27.600 12.900 30.000 22.500 ;
      LAYER met4 ;
        RECT 30.000 12.900 30.800 22.500 ;
      LAYER met4 ;
        RECT 30.800 12.900 33.200 22.500 ;
      LAYER met4 ;
        RECT 33.200 13.700 38.800 22.500 ;
        RECT 33.200 12.900 37.200 13.700 ;
      LAYER met4 ;
        RECT 37.200 12.900 38.000 13.700 ;
        RECT 22.000 12.100 29.200 12.900 ;
      LAYER met4 ;
        RECT 29.200 12.100 30.800 12.900 ;
      LAYER met4 ;
        RECT 30.800 12.100 34.800 12.900 ;
      LAYER met4 ;
        RECT 34.800 12.100 36.400 12.900 ;
      LAYER met4 ;
        RECT 36.400 12.100 38.000 12.900 ;
      LAYER met4 ;
        RECT 16.400 11.300 19.600 12.100 ;
      LAYER met4 ;
        RECT 19.600 11.300 20.400 12.100 ;
      LAYER met4 ;
        RECT 20.400 11.300 22.000 12.100 ;
      LAYER met4 ;
        RECT 22.000 11.300 28.400 12.100 ;
      LAYER met4 ;
        RECT 28.400 11.300 30.800 12.100 ;
      LAYER met4 ;
        RECT 30.800 11.300 38.000 12.100 ;
      LAYER met4 ;
        RECT 38.000 11.300 38.800 13.700 ;
      LAYER met4 ;
        RECT 38.800 12.900 41.200 22.500 ;
      LAYER met4 ;
        RECT 41.200 18.500 48.400 22.500 ;
      LAYER met4 ;
        RECT 48.400 18.500 50.800 22.500 ;
      LAYER met4 ;
        RECT 50.800 19.300 54.000 22.500 ;
      LAYER met4 ;
        RECT 54.000 20.900 56.400 22.500 ;
      LAYER met4 ;
        RECT 56.400 20.900 58.800 22.500 ;
      LAYER met4 ;
        RECT 54.000 20.100 55.600 20.900 ;
      LAYER met4 ;
        RECT 55.600 20.100 58.800 20.900 ;
      LAYER met4 ;
        RECT 54.000 19.300 54.800 20.100 ;
      LAYER met4 ;
        RECT 54.800 19.300 58.800 20.100 ;
        RECT 50.800 18.500 58.800 19.300 ;
      LAYER met4 ;
        RECT 58.800 18.500 61.200 22.500 ;
      LAYER met4 ;
        RECT 61.200 19.300 64.400 22.500 ;
      LAYER met4 ;
        RECT 64.400 20.900 66.800 22.500 ;
      LAYER met4 ;
        RECT 66.800 21.700 67.600 22.500 ;
      LAYER met4 ;
        RECT 67.600 21.700 75.600 22.500 ;
      LAYER met4 ;
        RECT 75.600 21.700 78.500 22.500 ;
        RECT 66.800 20.900 68.400 21.700 ;
      LAYER met4 ;
        RECT 68.400 20.900 76.400 21.700 ;
        RECT 64.400 20.100 66.000 20.900 ;
      LAYER met4 ;
        RECT 66.000 20.100 70.000 20.900 ;
      LAYER met4 ;
        RECT 70.000 20.100 76.400 20.900 ;
        RECT 64.400 19.300 65.200 20.100 ;
      LAYER met4 ;
        RECT 65.200 19.300 70.800 20.100 ;
        RECT 61.200 18.500 70.800 19.300 ;
        RECT 41.200 17.700 47.600 18.500 ;
      LAYER met4 ;
        RECT 47.600 17.700 53.200 18.500 ;
      LAYER met4 ;
        RECT 53.200 17.700 58.000 18.500 ;
      LAYER met4 ;
        RECT 58.000 17.700 63.600 18.500 ;
      LAYER met4 ;
        RECT 41.200 16.900 46.800 17.700 ;
      LAYER met4 ;
        RECT 46.800 16.900 53.200 17.700 ;
      LAYER met4 ;
        RECT 53.200 16.900 57.200 17.700 ;
      LAYER met4 ;
        RECT 57.200 16.900 63.600 17.700 ;
      LAYER met4 ;
        RECT 63.600 16.900 70.800 18.500 ;
        RECT 41.200 13.700 48.400 16.900 ;
        RECT 41.200 12.900 45.200 13.700 ;
      LAYER met4 ;
        RECT 45.200 12.900 46.000 13.700 ;
        RECT 38.800 12.100 42.800 12.900 ;
      LAYER met4 ;
        RECT 42.800 12.100 44.400 12.900 ;
      LAYER met4 ;
        RECT 44.400 12.100 46.000 12.900 ;
        RECT 38.800 11.300 46.000 12.100 ;
      LAYER met4 ;
        RECT 46.000 11.300 48.400 13.700 ;
      LAYER met4 ;
        RECT 48.400 11.300 50.800 16.900 ;
      LAYER met4 ;
        RECT 50.800 11.300 58.800 16.900 ;
      LAYER met4 ;
        RECT 58.800 12.900 61.200 16.900 ;
      LAYER met4 ;
        RECT 61.200 16.100 70.800 16.900 ;
        RECT 61.200 12.900 64.400 16.100 ;
      LAYER met4 ;
        RECT 64.400 15.300 65.200 16.100 ;
      LAYER met4 ;
        RECT 65.200 15.300 70.800 16.100 ;
      LAYER met4 ;
        RECT 64.400 14.500 66.000 15.300 ;
      LAYER met4 ;
        RECT 66.000 14.500 70.800 15.300 ;
      LAYER met4 ;
        RECT 64.400 12.900 66.800 14.500 ;
        RECT 58.800 11.300 66.800 12.900 ;
      LAYER met4 ;
        RECT 66.800 12.100 70.800 14.500 ;
      LAYER met4 ;
        RECT 70.800 12.900 73.200 20.100 ;
      LAYER met4 ;
        RECT 73.200 19.300 74.800 20.100 ;
      LAYER met4 ;
        RECT 74.800 19.300 76.400 20.100 ;
      LAYER met4 ;
        RECT 73.200 18.500 75.600 19.300 ;
      LAYER met4 ;
        RECT 75.600 18.500 76.400 19.300 ;
      LAYER met4 ;
        RECT 76.400 18.500 78.500 21.700 ;
        RECT 73.200 12.900 78.500 18.500 ;
      LAYER met4 ;
        RECT 70.800 12.100 74.800 12.900 ;
      LAYER met4 ;
        RECT 74.800 12.100 78.500 12.900 ;
        RECT 66.800 11.300 70.000 12.100 ;
      LAYER met4 ;
        RECT 70.000 11.300 74.000 12.100 ;
      LAYER met4 ;
        RECT 74.000 11.300 78.500 12.100 ;
        RECT 0.000 10.500 14.000 11.300 ;
      LAYER met4 ;
        RECT 14.000 10.500 14.800 11.300 ;
      LAYER met4 ;
        RECT 14.800 10.500 30.800 11.300 ;
      LAYER met4 ;
        RECT 30.800 10.500 31.600 11.300 ;
      LAYER met4 ;
        RECT 31.600 10.500 38.800 11.300 ;
      LAYER met4 ;
        RECT 38.800 10.500 39.600 11.300 ;
      LAYER met4 ;
        RECT 39.600 10.500 78.500 11.300 ;
        RECT 0.000 9.500 78.500 10.500 ;
  END
END qubitbytes_logo
END LIBRARY

