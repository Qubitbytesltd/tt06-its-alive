(* blackbox *)
module qubitbytes_logo_blackbox (
`ifdef USE_POWER_PINS
    input  VGND,
    input  VPWR
`endif  // USE_POWER_PINS
);
endmodule
