(* blackbox *)
module qubitbytes_logo (
`ifdef USE_POWER_PINS
    input  vss,
    input  vdd
`endif  // USE_POWER_PINS
);
endmodule
