  X �    ( �    (  skullfet_logo  >A�7KƧ�9D�/��ZT �    ( �    (  skullfet_logo     F   ,  ��      ��  � 2�  � 2�      ��          F   ,              �  ]�  �  ]�                  G   ,  P  [  P  ^$  -P  ^$  -P  [  P  [      G   ,  <�  [  <�  ^$  @  ^$  @  [  <�  [      G   ,  L�  [  L�  ^$  O�  ^$  O�  [  L�  [      G   ,  0  W�  0  [  -P  [  -P  W�  0  W�      G   ,  9�  W�  9�  [  @  [  @  W�  9�  W�      G   ,  Ip  W�  Ip  [  R�  [  R�  W�  Ip  W�      G   ,    E$    W�  p  W�  p  E$    E$      G   ,  #�  Q�  #�  W�  -P  W�  -P  Q�  #�  Q�      G   ,  #�  N�  #�  Q�  *0  Q�  *0  N�  #�  N�      G   ,  #�  Kd  #�  N�  '  N�  '  Kd  #�  Kd      G   ,  6�  Kd  6�  W�  @  W�  @  Kd  6�  Kd      G   ,  FP  T�  FP  W�  R�  W�  R�  T�  FP  T�      G   ,  C0  Q�  C0  T�  O�  T�  O�  Q�  C0  Q�      G   ,  C0  N�  C0  Q�  L�  Q�  L�  N�  C0  N�      G   ,  C0  Kd  C0  N�  Ip  N�  Ip  Kd  C0  Kd      G   ,  6�  HD  6�  Kd  Ip  Kd  Ip  HD  6�  HD      G   ,  3�  E$  3�  HD  FP  HD  FP  E$  3�  E$      G   ,  �  B  �  E$  -P  E$  -P  B  �  B      G   ,  0p  B  0p  E$  FP  E$  FP  B  0p  B      G   ,  
�  >�  
�  B  -P  B  -P  >�  
�  >�      G   ,  P  5�  P  8�  p  8�  p  5�  P  5�      G   ,  0  2d  0  5�  p  5�  p  2d  0  2d      G   ,  #�  2d  #�  >�  -P  >�  -P  2d  #�  2d      G   ,  6�  >�  6�  B  Ip  B  Ip  >�  6�  >�      G   ,    /D    2d  *0  2d  *0  /D    /D      G   ,  
�  ,$  
�  /D  '  /D  '  ,$  
�  ,$      G   ,  6�  ,$  6�  >�  @  >�  @  ,$  6�  ,$      G   ,  C0  ;�  C0  >�  Ip  >�  Ip  ;�  C0  ;�      G   ,  C0  8�  C0  ;�  L�  ;�  L�  8�  C0  8�      G   ,  C0  5�  C0  8�  O�  8�  O�  5�  C0  5�      G   ,  FP  2d  FP  5�  R�  5�  R�  2d  FP  2d      G   ,  Ip  /D  Ip  2d  R�  2d  R�  /D  Ip  /D      G   ,  U�  2d  U�  ^$  _P  ^$  _P  2d  U�  2d      G   ,  k�  [  k�  ^$  n�  ^$  n�  [  k�  [      G   ,  ~�  [  ~�  ^$  ��  ^$  ��  [  ~�  [      G   ,  ��  [  ��  ^$  ��  ^$  ��  [  ��  [      G   ,  �P  [  �P  ^$  �P  ^$  �P  [  �P  [      G   ,  ��  [  ��  ^$ �  ^$ �  [  ��  [      G   ,  k�  W�  k�  [  r  [  r  W�  k�  W�      G   ,  {p  W�  {p  [  ��  [  ��  W�  {p  W�      G   ,  ��  W�  ��  [  ��  [  ��  W�  ��  W�      G   ,  �0  W�  �0  [  �P  [  �P  W�  �0  W�      G   ,  ��  W�  ��  [ �  [ �  W�  ��  W�      G   , �  W� �  ^$ �  ^$ �  W� �  W�      G   ,  k�  2d  k�  W�  u0  W�  u0  2d  k�  2d      G   ,  xP  2d  xP  W�  ��  W�  ��  2d  xP  2d      G   ,  �P  2d  �P  5�  �p  5�  �p  2d  �P  2d      G   ,  U�  /D  U�  2d  r  2d  r  /D  U�  /D      G   ,  xP  /D  xP  2d  ��  2d  ��  /D  xP  /D      G   ,  �0  /D  �0  2d  �p  2d  �p  /D  �0  /D      G   ,  L�  ,$  L�  /D  O�  /D  O�  ,$  L�  ,$      G   ,  U�  ,$  U�  /D  n�  /D  n�  ,$  U�  ,$      G   ,  xP  ,$  xP  /D  �p  /D  �p  ,$  xP  ,$      G   ,  ��  2d  ��  W�  ��  W�  ��  2d  ��  2d      G   ,  �  HD  �  W�  �p  W�  �p  HD  �  HD      G   ,  ��  Q�  ��  W�  �P  W�  �P  Q�  ��  Q�      G   ,  ��  N�  ��  Q�  �0  Q�  �0  N�  ��  N�      G   ,  ��  Kd  ��  N�  �  N�  �  Kd  ��  Kd      G   ,  �  HD  �  W�  �  W�  �  HD  �  HD      G   ,  ��  Q�  ��  W� �  W� �  Q�  ��  Q�      G   ,   T�   W� 'P  W� 'P  T�   T�      G   , 0  Q� 0  T� *p  T� *p  Q� 0  Q�      G   ,  ��  N�  ��  Q� �  Q� �  N�  ��  N�      G   , p  N� p  Q� *p  Q� *p  N� p  N�      G   ,  ��  Kd  ��  N�  ��  N�  ��  Kd  ��  Kd      G   ,  ��  E$  ��  HD  ��  HD  ��  E$  ��  E$      G   ,  �  E$  �  HD  �p  HD  �p  E$  �  E$      G   ,  ��  B  ��  E$  ��  E$  ��  B  ��  B      G   ,  �p  B  �p  E$  �p  E$  �p  B  �p  B      G   ,  ��  2d  ��  5�  ��  5�  ��  2d  ��  2d      G   ,  ��  /D  ��  2d  �0  2d  �0  /D  ��  /D      G   ,  �p  /D  �p  2d  ��  2d  ��  /D  �p  /D      G   ,  ��  ,$  ��  /D  ��  /D  ��  ,$  ��  ,$      G   ,  �  ,$  �  B  �p  B  �p  ,$  �  ,$      G   ,  �  2d  �  B  �  B  �  2d  �  2d      G   ,  ��  ;�  ��  >�  ��  >�  ��  ;�  ��  ;�      G   ,  ��  8�  ��  ;� �  ;� �  8�  ��  8�      G   ,  ��  2d  ��  8� �  8� �  2d  ��  2d      G   ,  �  ,$  �  2d �  2d �  ,$  �  ,$      G   , �  2d �  N� �  N� �  2d �  2d      G   , $0  Kd $0  N� *p  N� *p  Kd $0  Kd      G   , 'P  HD 'P  Kd *p  Kd *p  HD 'P  HD      G   , �  /D �  2d $0  2d $0  /D �  /D      G   , p  ,$ p  /D !  /D !  ,$ p  ,$      G   ,  6�  )  6�  ,$  9�  ,$  9�  )  6�  )      G   ,  xP  )  xP  ,$  {p  ,$  {p  )  xP  )      G   ,  ��  )  ��  ,$  ��  ,$  ��  )  ��  )      F        @L������   .�  � VPWR      F        @L������  �  � VGND      F   ,  ��      ��  � 2�  � 2�      ��          F   ,              �  ]�  �  ]�                  H   ,  ��  jH  ��  k  �l  k  �l  jH  ��  jH      H   ,  �L  jH  �L  k  �  k  �  jH  �L  jH      H   ,  �l  jH  �l  k  �4  k  �4  jH  �l  jH      H   ,  �  jH  �  k  ��  k  ��  jH  �  jH      H   ,  ��  jH  ��  k  �L  k  �L  jH  ��  jH      H   ,  ��  jH  ��  k  ��  k  ��  jH  ��  jH      H   ,  ��  mh  ��  n0  �l  n0  �l  mh  ��  mh      H   ,  ��  l�  ��  mh  �l  mh  �l  l�  ��  l�      H   ,  ��  k�  ��  l�  �l  l�  �l  k�  ��  k�      H   ,  ��  k  ��  k�  �l  k�  �l  k  ��  k      H   ,  ��  r  ��  r�  �l  r�  �l  r  ��  r      H   ,  �L  v�  �L  w�  �  w�  �  v�  �L  v�      H   ,  �L  v   �L  v�  �  v�  �  v   �L  v       H   ,  �L  u8  �L  v   �  v   �  u8  �L  u8      H   ,  �L  tp  �L  u8  �  u8  �  tp  �L  tp      H   ,  �L  s�  �L  tp  �  tp  �  s�  �L  s�      H   ,  �L  r�  �L  s�  �  s�  �  r�  �L  r�      H   ,  �L  r  �L  r�  �  r�  �  r  �L  r      H   ,  �L  qP  �L  r  �  r  �  qP  �L  qP      H   ,  �L  p�  �L  qP  �  qP  �  p�  �L  p�      H   ,  �L  o�  �L  p�  �  p�  �  o�  �L  o�      H   ,  �L  n�  �L  o�  �  o�  �  n�  �L  n�      H   ,  �L  n0  �L  n�  �  n�  �  n0  �L  n0      H   ,  �L  mh  �L  n0  �  n0  �  mh  �L  mh      H   ,  �L  l�  �L  mh  �  mh  �  l�  �L  l�      H   ,  �L  k�  �L  l�  �  l�  �  k�  �L  k�      H   ,  �L  k  �L  k�  �  k�  �  k  �L  k      H   ,  ��  qP  ��  r  �l  r  �l  qP  ��  qP      H   ,  �l  o�  �l  p�  �4  p�  �4  o�  �l  o�      H   ,  �l  n�  �l  o�  �4  o�  �4  n�  �l  n�      H   ,  �l  n0  �l  n�  �4  n�  �4  n0  �l  n0      H   ,  �l  mh  �l  n0  �4  n0  �4  mh  �l  mh      H   ,  �l  l�  �l  mh  �4  mh  �4  l�  �l  l�      H   ,  �l  k�  �l  l�  �4  l�  �4  k�  �l  k�      H   ,  �l  k  �l  k�  �4  k�  �4  k  �l  k      H   ,  ��  p�  ��  qP  �l  qP  �l  p�  ��  p�      H   ,  ��  w�  ��  xX  ��  xX  ��  w�  ��  w�      H   ,  ��  v�  ��  w�  ��  w�  ��  v�  ��  v�      H   ,  ��  v   ��  v�  ��  v�  ��  v   ��  v       H   ,  ��  u8  ��  v   ��  v   ��  u8  ��  u8      H   ,  ��  tp  ��  u8  ��  u8  ��  tp  ��  tp      H   ,  ��  s�  ��  tp  ��  tp  ��  s�  ��  s�      H   ,  ��  r�  ��  s�  ��  s�  ��  r�  ��  r�      H   ,  ��  r  ��  r�  ��  r�  ��  r  ��  r      H   ,  ��  qP  ��  r  ��  r  ��  qP  ��  qP      H   ,  ��  p�  ��  qP  ��  qP  ��  p�  ��  p�      H   ,  �  v   �  v�  ��  v�  ��  v   �  v       H   ,  �  u8  �  v   ��  v   ��  u8  �  u8      H   ,  �  tp  �  u8  ��  u8  ��  tp  �  tp      H   ,  �  s�  �  tp  ��  tp  ��  s�  �  s�      H   ,  �  r�  �  s�  ��  s�  ��  r�  �  r�      H   ,  �  r  �  r�  ��  r�  ��  r  �  r      H   ,  �  qP  �  r  ��  r  ��  qP  �  qP      H   ,  �  p�  �  qP  ��  qP  ��  p�  �  p�      H   ,  �  o�  �  p�  ��  p�  ��  o�  �  o�      H   ,  �  n�  �  o�  ��  o�  ��  n�  �  n�      H   ,  �  n0  �  n�  ��  n�  ��  n0  �  n0      H   ,  �  mh  �  n0  ��  n0  ��  mh  �  mh      H   ,  �  l�  �  mh  ��  mh  ��  l�  �  l�      H   ,  �  k�  �  l�  ��  l�  ��  k�  �  k�      H   ,  �  k  �  k�  ��  k�  ��  k  �  k      H   ,  ��  o�  ��  p�  �l  p�  �l  o�  ��  o�      H   ,  ��  v�  ��  w�  �L  w�  �L  v�  ��  v�      H   ,  ��  v   ��  v�  �L  v�  �L  v   ��  v       H   ,  ��  u8  ��  v   �L  v   �L  u8  ��  u8      H   ,  ��  tp  ��  u8  �L  u8  �L  tp  ��  tp      H   ,  ��  s�  ��  tp  �L  tp  �L  s�  ��  s�      H   ,  ��  r�  ��  s�  �L  s�  �L  r�  ��  r�      H   ,  ��  r  ��  r�  �L  r�  �L  r  ��  r      H   ,  ��  qP  ��  r  �L  r  �L  qP  ��  qP      H   ,  ��  p�  ��  qP  �L  qP  �L  p�  ��  p�      H   ,  ��  o�  ��  p�  �L  p�  �L  o�  ��  o�      H   ,  ��  n�  ��  o�  �L  o�  �L  n�  ��  n�      H   ,  ��  n0  ��  n�  �L  n�  �L  n0  ��  n0      H   ,  ��  mh  ��  n0  �L  n0  �L  mh  ��  mh      H   ,  ��  l�  ��  mh  �L  mh  �L  l�  ��  l�      H   ,  ��  k�  ��  l�  �L  l�  �L  k�  ��  k�      H   ,  ��  tp  ��  u8  ��  u8  ��  tp  ��  tp      H   ,  ��  k  ��  k�  �L  k�  �L  k  ��  k      H   ,  ��  s�  ��  tp  ��  tp  ��  s�  ��  s�      H   ,  ��  n�  ��  o�  �l  o�  �l  n�  ��  n�      H   ,  ��  r�  ��  s�  ��  s�  ��  r�  ��  r�      H   ,  ��  r  ��  r�  ��  r�  ��  r  ��  r      H   ,  ��  qP  ��  r  ��  r  ��  qP  ��  qP      H   ,  ��  p�  ��  qP  ��  qP  ��  p�  ��  p�      H   ,  ��  o�  ��  p�  ��  p�  ��  o�  ��  o�      H   ,  ��  n�  ��  o�  ��  o�  ��  n�  ��  n�      H   ,  ��  n0  ��  n�  ��  n�  ��  n0  ��  n0      H   ,  ��  mh  ��  n0  ��  n0  ��  mh  ��  mh      H   ,  ��  l�  ��  mh  ��  mh  ��  l�  ��  l�      H   ,  ��  k�  ��  l�  ��  l�  ��  k�  ��  k�      H   ,  ��  k  ��  k�  ��  k�  ��  k  ��  k      H   ,  ��  n0  ��  n�  �l  n�  �l  n0  ��  n0      H   ,  ��  r�  ��  s�  �l  s�  �l  r�  ��  r�      H   ,  ��  ]   ��  ]�  ��  ]�  ��  ]   ��  ]       H   ,  �L  `   �L  `�  �  `�  �  `   �L  `       H   ,  �L  _X  �L  `   �  `   �  _X  �L  _X      H   ,  �L  ^�  �L  _X  �  _X  �  ^�  �L  ^�      H   ,  �L  ]�  �L  ^�  �  ^�  �  ]�  �L  ]�      H   ,  �L  ]   �L  ]�  �  ]�  �  ]   �L  ]       H   ,  ��  g�  ��  h�  �l  h�  �l  g�  ��  g�      H   ,  ��  a�  ��  bx  �l  bx  �l  a�  ��  a�      H   ,  ��  e�  ��  f`  �l  f`  �l  e�  ��  e�      H   ,  ��  i�  ��  jH  �l  jH  �l  i�  ��  i�      H   ,  ��  d�  ��  e�  �l  e�  �l  d�  ��  d�      H   ,  ��  g(  ��  g�  �l  g�  �l  g(  ��  g(      H   ,  �  i�  �  jH  ��  jH  ��  i�  �  i�      H   ,  �  h�  �  i�  ��  i�  ��  h�  �  h�      H   ,  �  g�  �  h�  ��  h�  ��  g�  �  g�      H   ,  �  g(  �  g�  ��  g�  ��  g(  �  g(      H   ,  �  f`  �  g(  ��  g(  ��  f`  �  f`      H   ,  �  e�  �  f`  ��  f`  ��  e�  �  e�      H   ,  �  d�  �  e�  ��  e�  ��  d�  �  d�      H   ,  �  d  �  d�  ��  d�  ��  d  �  d      H   ,  �  c@  �  d  ��  d  ��  c@  �  c@      H   ,  �  bx  �  c@  ��  c@  ��  bx  �  bx      H   ,  �  a�  �  bx  ��  bx  ��  a�  �  a�      H   ,  �  `�  �  a�  ��  a�  ��  `�  �  `�      H   ,  �  `   �  `�  ��  `�  ��  `   �  `       H   ,  �  _X  �  `   ��  `   ��  _X  �  _X      H   ,  �  ^�  �  _X  ��  _X  ��  ^�  �  ^�      H   ,  �  ]�  �  ^�  ��  ^�  ��  ]�  �  ]�      H   ,  �  ]   �  ]�  ��  ]�  ��  ]   �  ]       H   ,  ��  d  ��  d�  �l  d�  �l  d  ��  d      H   ,  ��  h�  ��  i�  �l  i�  �l  h�  ��  h�      H   ,  �l  i�  �l  jH  �4  jH  �4  i�  �l  i�      H   ,  �l  h�  �l  i�  �4  i�  �4  h�  �l  h�      H   ,  �l  g�  �l  h�  �4  h�  �4  g�  �l  g�      H   ,  �l  g(  �l  g�  �4  g�  �4  g(  �l  g(      H   ,  ��  c@  ��  d  �l  d  �l  c@  ��  c@      H   ,  ��  f`  ��  g(  �l  g(  �l  f`  ��  f`      H   ,  ��  bx  ��  c@  �l  c@  �l  bx  ��  bx      H   ,  �L  i�  �L  jH  �  jH  �  i�  �L  i�      H   ,  �L  h�  �L  i�  �  i�  �  h�  �L  h�      H   ,  �L  g�  �L  h�  �  h�  �  g�  �L  g�      H   ,  �L  g(  �L  g�  �  g�  �  g(  �L  g(      H   ,  �L  f`  �L  g(  �  g(  �  f`  �L  f`      H   ,  �L  e�  �L  f`  �  f`  �  e�  �L  e�      H   ,  �L  d�  �L  e�  �  e�  �  d�  �L  d�      H   ,  ��  e�  ��  f`  ��  f`  ��  e�  ��  e�      H   ,  ��  d�  ��  e�  ��  e�  ��  d�  ��  d�      H   ,  ��  d  ��  d�  ��  d�  ��  d  ��  d      H   ,  ��  c@  ��  d  ��  d  ��  c@  ��  c@      H   ,  ��  i�  ��  jH  �L  jH  �L  i�  ��  i�      H   ,  ��  bx  ��  c@  ��  c@  ��  bx  ��  bx      H   ,  ��  h�  ��  i�  �L  i�  �L  h�  ��  h�      H   ,  ��  a�  ��  bx  ��  bx  ��  a�  ��  a�      H   ,  ��  g�  ��  h�  �L  h�  �L  g�  ��  g�      H   ,  ��  `�  ��  a�  ��  a�  ��  `�  ��  `�      H   ,  ��  g(  ��  g�  �L  g�  �L  g(  ��  g(      H   ,  �L  d  �L  d�  �  d�  �  d  �L  d      H   ,  ��  f`  ��  g(  �L  g(  �L  f`  ��  f`      H   ,  ��  `   ��  `�  ��  `�  ��  `   ��  `       H   ,  ��  e�  ��  f`  �L  f`  �L  e�  ��  e�      H   ,  �L  c@  �L  d  �  d  �  c@  �L  c@      H   ,  ��  d�  ��  e�  �L  e�  �L  d�  ��  d�      H   ,  ��  _X  ��  `   ��  `   ��  _X  ��  _X      H   ,  ��  d  ��  d�  �L  d�  �L  d  ��  d      H   ,  �L  bx  �L  c@  �  c@  �  bx  �L  bx      H   ,  ��  c@  ��  d  �L  d  �L  c@  ��  c@      H   ,  ��  ^�  ��  _X  ��  _X  ��  ^�  ��  ^�      H   ,  ��  bx  ��  c@  �L  c@  �L  bx  ��  bx      H   ,  �L  a�  �L  bx  �  bx  �  a�  �L  a�      H   ,  ��  a�  ��  bx  �L  bx  �L  a�  ��  a�      H   ,  ��  ]�  ��  ^�  ��  ^�  ��  ]�  ��  ]�      H   ,  ��  `�  ��  a�  �L  a�  �L  `�  ��  `�      H   ,  ��  i�  ��  jH  ��  jH  ��  i�  ��  i�      H   ,  ��  `   ��  `�  �L  `�  �L  `   ��  `       H   ,  ��  h�  ��  i�  ��  i�  ��  h�  ��  h�      H   ,  ��  _X  ��  `   �L  `   �L  _X  ��  _X      H   ,  ��  g�  ��  h�  ��  h�  ��  g�  ��  g�      H   ,  ��  ^�  ��  _X  �L  _X  �L  ^�  ��  ^�      H   ,  ��  g(  ��  g�  ��  g�  ��  g(  ��  g(      H   ,  ��  ]�  ��  ^�  �L  ^�  �L  ]�  ��  ]�      H   ,  ��  f`  ��  g(  ��  g(  ��  f`  ��  f`      H   ,  ��  ]   ��  ]�  �L  ]�  �L  ]   ��  ]       H   ,  ��  e�  ��  f`  ��  f`  ��  e�  ��  e�      H   ,  ��  d�  ��  e�  ��  e�  ��  d�  ��  d�      H   ,  ��  d  ��  d�  ��  d�  ��  d  ��  d      H   ,  ��  c@  ��  d  ��  d  ��  c@  ��  c@      H   ,  ��  bx  ��  c@  ��  c@  ��  bx  ��  bx      H   ,  ��  a�  ��  bx  ��  bx  ��  a�  ��  a�      H   ,  ��  `�  ��  a�  ��  a�  ��  `�  ��  `�      H   ,  ��  `   ��  `�  ��  `�  ��  `   ��  `       H   ,  ��  _X  ��  `   ��  `   ��  _X  ��  _X      H   ,  ��  ^�  ��  _X  ��  _X  ��  ^�  ��  ^�      H   ,  ��  ]�  ��  ^�  ��  ^�  ��  ]�  ��  ]�      H   ,  �L  `�  �L  a�  �  a�  �  `�  �L  `�      H   ,  �4  jH  �4  k  ��  k  ��  jH  �4  jH      H   ,  �T  jH  �T  k  �  k  �  jH  �T  jH      H   ,  ��  jH  ��  k  ��  k  ��  jH  ��  jH      H   ,  ��  r  ��  r�  �t  r�  �t  r  ��  r      H   ,  ��  qP  ��  r  �t  r  �t  qP  ��  qP      H   ,  ��  p�  ��  qP  �t  qP  �t  p�  ��  p�      H   ,  ��  o�  ��  p�  �t  p�  �t  o�  ��  o�      H   ,  ��  n�  ��  o�  �t  o�  �t  n�  ��  n�      H   ,  �l  jH  �l  k  �4  k  �4  jH  �l  jH      H   ,  ��  n0  ��  n�  �t  n�  �t  n0  ��  n0      H   ,  ��  mh  ��  n0  �t  n0  �t  mh  ��  mh      H   ,  ��  l�  ��  mh  �t  mh  �t  l�  ��  l�      H   ,  ��  k�  ��  l�  �t  l�  �t  k�  ��  k�      H   ,  ��  jH  ��  k  ��  k  ��  jH  ��  jH      H   ,  ��  jH  ��  k  ��  k  ��  jH  ��  jH      H   ,  �  jH  �  k  ��  k  ��  jH  �  jH      H   ,  ��  jH  ��  k  �T  k  �T  jH  ��  jH      H   ,  ��  jH  ��  k  �l  k  �l  jH  ��  jH      H   ,  ��  u8  ��  v   �|  v   �|  u8  ��  u8      H   ,  ��  tp  ��  u8  �|  u8  �|  tp  ��  tp      H   ,  ��  s�  ��  tp  �|  tp  �|  s�  ��  s�      H   ,  ��  r�  ��  s�  �|  s�  �|  r�  ��  r�      H   ,  ��  r  ��  r�  �|  r�  �|  r  ��  r      H   ,  ��  qP  ��  r  ��  r  ��  qP  ��  qP      H   ,  ��  qP  ��  r  �\  r  �\  qP  ��  qP      H   ,  �$  qP  �$  r  ��  r  ��  qP  �$  qP      H   ,  �<  qP  �<  r  �  r  �  qP  �<  qP      H   ,  ��  qP  ��  r  ��  r  ��  qP  ��  qP      H   ,  ��  v�  ��  w�  �|  w�  �|  v�  ��  v�      H   ,  �  qP  �  r  ��  r  ��  qP  �  qP      H   ,  �t  qP  �t  r  �<  r  �<  qP  �t  qP      H   ,  �\  qP  �\  r  �$  r  �$  qP  �\  qP      H   ,  ��  v   ��  v�  �|  v�  �|  v   ��  v       H   ,  �d  w�  �d  xX  �,  xX  �,  w�  �d  w�      H   ,  �d  v�  �d  w�  �,  w�  �,  v�  �d  v�      H   ,  �  u8  �  v   ��  v   ��  u8  �  u8      H   ,  �d  v   �d  v�  �,  v�  �,  v   �d  v       H   ,  ��  r�  ��  s�  ��  s�  ��  r�  ��  r�      H   ,  �d  u8  �d  v   �,  v   �,  u8  �d  u8      H   ,  �d  tp  �d  u8  �,  u8  �,  tp  �d  tp      H   ,  �  tp  �  u8  ��  u8  ��  tp  �  tp      H   ,  �d  s�  �d  tp  �,  tp  �,  s�  �d  s�      H   ,  ��  r  ��  r�  ��  r�  ��  r  ��  r      H   ,  �  s�  �  tp  ��  tp  ��  s�  �  s�      H   ,  �|  w�  �|  xX  �D  xX  �D  w�  �|  w�      H   ,  �|  v�  �|  w�  �D  w�  �D  v�  �|  v�      H   ,  �|  v   �|  v�  �D  v�  �D  v   �|  v       H   ,  �|  u8  �|  v   �D  v   �D  u8  �|  u8      H   ,  �|  tp  �|  u8  �D  u8  �D  tp  �|  tp      H   ,  �|  s�  �|  tp  �D  tp  �D  s�  �|  s�      H   ,  �|  r�  �|  s�  �D  s�  �D  r�  �|  r�      H   ,  ��  u8  ��  v   �d  v   �d  u8  ��  u8      H   ,  ��  w�  ��  xX  �d  xX  �d  w�  ��  w�      H   ,  ��  v�  ��  w�  ��  w�  ��  v�  ��  v�      H   ,  ��  tp  ��  u8  �d  u8  �d  tp  ��  tp      H   ,  ��  v   ��  v�  ��  v�  ��  v   ��  v       H   ,  �  w�  �  xX  ��  xX  ��  w�  �  w�      H   ,  ��  u8  ��  v   ��  v   ��  u8  ��  u8      H   ,  ��  w�  ��  xX  ��  xX  ��  w�  ��  w�      H   ,  ��  v   ��  v�  �d  v�  �d  v   ��  v       H   ,  ��  v�  ��  w�  ��  w�  ��  v�  ��  v�      H   ,  ��  v   ��  v�  ��  v�  ��  v   ��  v       H   ,  ��  u8  ��  v   ��  v   ��  u8  ��  u8      H   ,  ��  s�  ��  tp  �d  tp  �d  s�  ��  s�      H   ,  ��  tp  ��  u8  ��  u8  ��  tp  ��  tp      H   ,  ��  s�  ��  tp  ��  tp  ��  s�  ��  s�      H   ,  ��  w�  ��  xX  ��  xX  ��  w�  ��  w�      H   ,  �  v�  �  w�  ��  w�  ��  v�  �  v�      H   ,  ��  tp  ��  u8  ��  u8  ��  tp  ��  tp      H   ,  �,  w�  �,  xX  ��  xX  ��  w�  �,  w�      H   ,  �,  v�  �,  w�  ��  w�  ��  v�  �,  v�      H   ,  ��  v�  ��  w�  �d  w�  �d  v�  ��  v�      H   ,  �,  v   �,  v�  ��  v�  ��  v   �,  v       H   ,  �,  u8  �,  v   ��  v   ��  u8  �,  u8      H   ,  �,  tp  �,  u8  ��  u8  ��  tp  �,  tp      H   ,  �,  s�  �,  tp  ��  tp  ��  s�  �,  s�      H   ,  �D  w�  �D  xX  �  xX  �  w�  �D  w�      H   ,  �  v   �  v�  ��  v�  ��  v   �  v       H   ,  �D  v�  �D  w�  �  w�  �  v�  �D  v�      H   ,  �D  v   �D  v�  �  v�  �  v   �D  v       H   ,  �D  u8  �D  v   �  v   �  u8  �D  u8      H   ,  �D  tp  �D  u8  �  u8  �  tp  �D  tp      H   ,  �D  s�  �D  tp  �  tp  �  s�  �D  s�      H   ,  �D  r�  �D  s�  �  s�  �  r�  �D  r�      H   ,  ��  s�  ��  tp  ��  tp  ��  s�  ��  s�      H   ,  ��  s�  ��  tp  �\  tp  �\  s�  ��  s�      H   ,  �$  s�  �$  tp  ��  tp  ��  s�  �$  s�      H   ,  �$  r  �$  r�  ��  r�  ��  r  �$  r      H   ,  �  tp  �  u8  ��  u8  ��  tp  �  tp      H   ,  ��  r�  ��  s�  �\  s�  �\  r�  ��  r�      H   ,  �  s�  �  tp  ��  tp  ��  s�  �  s�      H   ,  ��  r  ��  r�  �\  r�  �\  r  ��  r      H   ,  �  r�  �  s�  ��  s�  ��  r�  �  r�      H   ,  �  r  �  r�  ��  r�  ��  r  �  r      H   ,  �$  r�  �$  s�  ��  s�  ��  r�  �$  r�      H   ,  �$  v   �$  v�  ��  v�  ��  v   �$  v       H   ,  ��  u8  ��  v   ��  v   ��  u8  ��  u8      H   ,  ��  tp  ��  u8  ��  u8  ��  tp  ��  tp      H   ,  �t  r�  �t  s�  �<  s�  �<  r�  �t  r�      H   ,  ��  s�  ��  tp  ��  tp  ��  s�  ��  s�      H   ,  �t  r  �t  r�  �<  r�  �<  r  �t  r      H   ,  ��  r�  ��  s�  ��  s�  ��  r�  ��  r�      H   ,  ��  v�  ��  w�  ��  w�  ��  v�  ��  v�      H   ,  �$  tp  �$  u8  ��  u8  ��  tp  �$  tp      H   ,  ��  v   ��  v�  ��  v�  ��  v   ��  v       H   ,  ��  u8  ��  v   ��  v   ��  u8  ��  u8      H   ,  �\  v   �\  v�  �$  v�  �$  v   �\  v       H   ,  ��  r  ��  r�  ��  r�  ��  r  ��  r      H   ,  �\  u8  �\  v   �$  v   �$  u8  �\  u8      H   ,  �\  tp  �\  u8  �$  u8  �$  tp  �\  tp      H   ,  �\  s�  �\  tp  �$  tp  �$  s�  �\  s�      H   ,  �\  r�  �\  s�  �$  s�  �$  r�  �\  r�      H   ,  �\  r  �\  r�  �$  r�  �$  r  �\  r      H   ,  ��  tp  ��  u8  ��  u8  ��  tp  ��  tp      H   ,  �<  r�  �<  s�  �  s�  �  r�  �<  r�      H   ,  ��  s�  ��  tp  ��  tp  ��  s�  ��  s�      H   ,  ��  r�  ��  s�  ��  s�  ��  r�  ��  r�      H   ,  ��  r  ��  r�  ��  r�  ��  r  ��  r      H   ,  ��  u8  ��  v   �\  v   �\  u8  ��  u8      H   ,  �<  s�  �<  tp  �  tp  �  s�  �<  s�      H   ,  �$  u8  �$  v   ��  v   ��  u8  �$  u8      H   ,  ��  tp  ��  u8  �\  u8  �\  tp  ��  tp      H   ,  �<  r  �<  r�  �  r�  �  r  �<  r      H   ,  �  n�  �  o�  ��  o�  ��  n�  �  n�      H   ,  �  n0  �  n�  ��  n�  ��  n0  �  n0      H   ,  �t  n0  �t  n�  �<  n�  �<  n0  �t  n0      H   ,  ��  n�  ��  o�  ��  o�  ��  n�  ��  n�      H   ,  �t  mh  �t  n0  �<  n0  �<  mh  �t  mh      H   ,  �<  o�  �<  p�  �  p�  �  o�  �<  o�      H   ,  �t  l�  �t  mh  �<  mh  �<  l�  �t  l�      H   ,  �<  n0  �<  n�  �  n�  �  n0  �<  n0      H   ,  ��  o�  ��  p�  ��  p�  ��  o�  ��  o�      H   ,  �<  mh  �<  n0  �  n0  �  mh  �<  mh      H   ,  ��  p�  ��  qP  �\  qP  �\  p�  ��  p�      H   ,  �<  p�  �<  qP  �  qP  �  p�  �<  p�      H   ,  ��  p�  ��  qP  ��  qP  ��  p�  ��  p�      H   ,  �\  p�  �\  qP  �$  qP  �$  p�  �\  p�      H   ,  �<  n�  �<  o�  �  o�  �  n�  �<  n�      H   ,  ��  o�  ��  p�  �\  p�  �\  o�  ��  o�      H   ,  �t  p�  �t  qP  �<  qP  �<  p�  �t  p�      H   ,  �  p�  �  qP  ��  qP  ��  p�  �  p�      H   ,  �t  o�  �t  p�  �<  p�  �<  o�  �t  o�      H   ,  �  o�  �  p�  ��  p�  ��  o�  �  o�      H   ,  �t  n�  �t  o�  �<  o�  �<  n�  �t  n�      H   ,  ��  k  ��  k�  ��  k�  ��  k  ��  k      H   ,  �T  k�  �T  l�  �  l�  �  k�  �T  k�      H   ,  ��  mh  ��  n0  ��  n0  ��  mh  ��  mh      H   ,  ��  l�  ��  mh  ��  mh  ��  l�  ��  l�      H   ,  �  p�  �  qP  ��  qP  ��  p�  �  p�      H   ,  �4  l�  �4  mh  ��  mh  ��  l�  �4  l�      H   ,  ��  k�  ��  l�  ��  l�  ��  k�  ��  k�      H   ,  ��  k  ��  k�  ��  k�  ��  k  ��  k      H   ,  �  o�  �  p�  ��  p�  ��  o�  �  o�      H   ,  �T  o�  �T  p�  �  p�  �  o�  �T  o�      H   ,  ��  o�  ��  p�  ��  p�  ��  o�  ��  o�      H   ,  �  n�  �  o�  ��  o�  ��  n�  �  n�      H   ,  ��  mh  ��  n0  ��  n0  ��  mh  ��  mh      H   ,  �  n0  �  n�  ��  n�  ��  n0  �  n0      H   ,  �4  k�  �4  l�  ��  l�  ��  k�  �4  k�      H   ,  �  mh  �  n0  ��  n0  ��  mh  �  mh      H   ,  �T  k  �T  k�  �  k�  �  k  �T  k      H   ,  ��  l�  ��  mh  ��  mh  ��  l�  ��  l�      H   ,  �  l�  �  mh  ��  mh  ��  l�  �  l�      H   ,  ��  n�  ��  o�  ��  o�  ��  n�  ��  n�      H   ,  �4  k  �4  k�  ��  k�  ��  k  �4  k      H   ,  �  k�  �  l�  ��  l�  ��  k�  �  k�      H   ,  �l  k�  �l  l�  �4  l�  �4  k�  �l  k�      H   ,  �  k  �  k�  ��  k�  ��  k  �  k      H   ,  ��  n0  ��  n�  ��  n�  ��  n0  ��  n0      H   ,  ��  n�  ��  o�  �T  o�  �T  n�  ��  n�      H   ,  �T  n�  �T  o�  �  o�  �  n�  �T  n�      H   ,  ��  n0  ��  n�  �T  n�  �T  n0  ��  n0      H   ,  �T  n0  �T  n�  �  n�  �  n0  �T  n0      H   ,  ��  k�  ��  l�  ��  l�  ��  k�  ��  k�      H   ,  ��  mh  ��  n0  �T  n0  �T  mh  ��  mh      H   ,  ��  mh  ��  n0  ��  n0  ��  mh  ��  mh      H   ,  ��  qP  ��  r  ��  r  ��  qP  ��  qP      H   ,  ��  l�  ��  mh  �T  mh  �T  l�  ��  l�      H   ,  ��  l�  ��  mh  ��  mh  ��  l�  ��  l�      H   ,  �T  mh  �T  n0  �  n0  �  mh  �T  mh      H   ,  ��  k�  ��  l�  �T  l�  �T  k�  ��  k�      H   ,  �l  k  �l  k�  �4  k�  �4  k  �l  k      H   ,  ��  k  ��  k�  �T  k�  �T  k  ��  k      H   ,  ��  k�  ��  l�  ��  l�  ��  k�  ��  k�      H   ,  ��  p�  ��  qP  ��  qP  ��  p�  ��  p�      H   ,  ��  k  ��  k�  ��  k�  ��  k  ��  k      H   ,  ��  n0  ��  n�  ��  n�  ��  n0  ��  n0      H   ,  ��  k  ��  k�  �l  k�  �l  k  ��  k      H   ,  �T  l�  �T  mh  �  mh  �  l�  �T  l�      H   ,  �  c@  �  d  ��  d  ��  c@  �  c@      H   ,  ��  c@  ��  d  �l  d  �l  c@  ��  c@      H   ,  �,  c@  �,  d  ��  d  ��  c@  �,  c@      H   ,  ��  g(  ��  g�  �l  g�  �l  g(  ��  g(      H   ,  �L  c@  �L  d  �  d  �  c@  �L  c@      H   ,  ��  c@  ��  d  �L  d  �L  c@  ��  c@      H   ,  ��  c@  ��  d  ��  d  ��  c@  ��  c@      H   ,  ��  c@  ��  d  ��  d  ��  c@  ��  c@      H   ,  ��  h�  ��  i�  �l  i�  �l  h�  ��  h�      H   ,  ��  e�  ��  f`  �l  f`  �l  e�  ��  e�      H   ,  ��  g�  ��  h�  �l  h�  �l  g�  ��  g�      H   ,  ��  f`  ��  g(  �l  g(  �l  f`  ��  f`      H   ,  ��  d  ��  d�  �l  d�  �l  d  ��  d      H   ,  ��  c@  ��  d  ��  d  ��  c@  ��  c@      H   ,  ��  i�  ��  jH  �l  jH  �l  i�  ��  i�      H   ,  ��  d�  ��  e�  �l  e�  �l  d�  ��  d�      H   ,  ��  f`  ��  g(  ��  g(  ��  f`  ��  f`      H   ,  �l  i�  �l  jH  �4  jH  �4  i�  �l  i�      H   ,  ��  h�  ��  i�  ��  i�  ��  h�  ��  h�      H   ,  ��  g�  ��  h�  ��  h�  ��  g�  ��  g�      H   ,  �l  h�  �l  i�  �4  i�  �4  h�  �l  h�      H   ,  �4  e�  �4  f`  ��  f`  ��  e�  �4  e�      H   ,  �l  g�  �l  h�  �4  h�  �4  g�  �l  g�      H   ,  �l  g(  �l  g�  �4  g�  �4  g(  �l  g(      H   ,  �l  f`  �l  g(  �4  g(  �4  f`  �l  f`      H   ,  �T  i�  �T  jH  �  jH  �  i�  �T  i�      H   ,  �l  e�  �l  f`  �4  f`  �4  e�  �l  e�      H   ,  �l  d�  �l  e�  �4  e�  �4  d�  �l  d�      H   ,  �4  h�  �4  i�  ��  i�  ��  h�  �4  h�      H   ,  ��  i�  ��  jH  ��  jH  ��  i�  ��  i�      H   ,  ��  h�  ��  i�  ��  i�  ��  h�  ��  h�      H   ,  ��  g�  ��  h�  ��  h�  ��  g�  ��  g�      H   ,  ��  g(  ��  g�  ��  g�  ��  g(  ��  g(      H   ,  �4  g�  �4  h�  ��  h�  ��  g�  �4  g�      H   ,  ��  i�  ��  jH  �T  jH  �T  i�  ��  i�      H   ,  ��  h�  ��  i�  �T  i�  �T  h�  ��  h�      H   ,  �4  g(  �4  g�  ��  g�  ��  g(  �4  g(      H   ,  ��  i�  ��  jH  ��  jH  ��  i�  ��  i�      H   ,  �4  f`  �4  g(  ��  g(  ��  f`  �4  f`      H   ,  �4  i�  �4  jH  ��  jH  ��  i�  �4  i�      H   ,  �  f`  �  g(  ��  g(  ��  f`  �  f`      H   ,  �  e�  �  f`  ��  f`  ��  e�  �  e�      H   ,  �L  f`  �L  g(  �  g(  �  f`  �L  f`      H   ,  ��  e�  ��  f`  �L  f`  �L  e�  ��  e�      H   ,  �  d�  �  e�  ��  e�  ��  d�  �  d�      H   ,  �L  g�  �L  h�  �  h�  �  g�  �L  g�      H   ,  �  d  �  d�  ��  d�  ��  d  �  d      H   ,  �L  e�  �L  f`  �  f`  �  e�  �L  e�      H   ,  ��  i�  ��  jH  ��  jH  ��  i�  ��  i�      H   ,  ��  g(  ��  g�  �L  g�  �L  g(  ��  g(      H   ,  ��  d�  ��  e�  �L  e�  �L  d�  ��  d�      H   ,  ��  h�  ��  i�  ��  i�  ��  h�  ��  h�      H   ,  �  g�  �  h�  ��  h�  ��  g�  �  g�      H   ,  ��  g�  ��  h�  ��  h�  ��  g�  ��  g�      H   ,  �  g(  �  g�  ��  g�  ��  g(  �  g(      H   ,  ��  g(  ��  g�  ��  g�  ��  g(  ��  g(      H   ,  ��  f`  ��  g(  �L  g(  �L  f`  ��  f`      H   ,  �L  d�  �L  e�  �  e�  �  d�  �L  d�      H   ,  ��  d  ��  d�  �L  d�  �L  d  ��  d      H   ,  ��  f`  ��  g(  ��  g(  ��  f`  ��  f`      H   ,  ��  d�  ��  e�  ��  e�  ��  d�  ��  d�      H   ,  ��  e�  ��  f`  ��  f`  ��  e�  ��  e�      H   ,  �L  d  �L  d�  �  d�  �  d  �L  d      H   ,  ��  e�  ��  f`  ��  f`  ��  e�  ��  e�      H   ,  ��  d�  ��  e�  ��  e�  ��  d�  ��  d�      H   ,  ��  d  ��  d�  ��  d�  ��  d  ��  d      H   ,  ��  d  ��  d�  ��  d�  ��  d  ��  d      H   ,  ��  d�  ��  e�  ��  e�  ��  d�  ��  d�      H   ,  �L  g(  �L  g�  �  g�  �  g(  �L  g(      H   ,  �  h�  �  i�  ��  i�  ��  h�  �  h�      H   ,  ��  d  ��  d�  ��  d�  ��  d  ��  d      H   ,  ��  `   ��  `�  ��  `�  ��  `   ��  `       H   ,  ��  `�  ��  a�  ��  a�  ��  `�  ��  `�      H   ,  �d  `�  �d  a�  �,  a�  �,  `�  �d  `�      H   ,  ��  `�  ��  a�  �L  a�  �L  `�  ��  `�      H   ,  �,  a�  �,  bx  ��  bx  ��  a�  �,  a�      H   ,  �L  a�  �L  bx  �  bx  �  a�  �L  a�      H   ,  �  bx  �  c@  ��  c@  ��  bx  �  bx      H   ,  �d  `   �d  `�  �,  `�  �,  `   �d  `       H   ,  �  a�  �  bx  ��  bx  ��  a�  �  a�      H   ,  ��  `   ��  `�  �L  `�  �L  `   ��  `       H   ,  �L  `�  �L  a�  �  a�  �  `�  �L  `�      H   ,  �d  _X  �d  `   �,  `   �,  _X  �d  _X      H   ,  �,  _X  �,  `   ��  `   ��  _X  �,  _X      H   ,  �,  `   �,  `�  ��  `�  ��  `   �,  `       H   ,  ��  _X  ��  `   �L  `   �L  _X  ��  _X      H   ,  �,  bx  �,  c@  ��  c@  ��  bx  �,  bx      H   ,  �L  bx  �L  c@  �  c@  �  bx  �L  bx      H   ,  �d  ^�  �d  _X  �,  _X  �,  ^�  �d  ^�      H   ,  ��  bx  ��  c@  ��  c@  ��  bx  ��  bx      H   ,  ��  a�  ��  bx  ��  bx  ��  a�  ��  a�      H   ,  ��  _X  ��  `   ��  `   ��  _X  ��  _X      H   ,  �d  ]�  �d  ^�  �,  ^�  �,  ]�  �d  ]�      H   ,  �L  `   �L  `�  �  `�  �  `   �L  `       H   ,  ��  bx  ��  c@  �L  c@  �L  bx  ��  bx      H   ,  �d  ]   �d  ]�  �,  ]�  �,  ]   �d  ]       H   ,  ��  a�  ��  bx  ��  bx  ��  a�  ��  a�      H   ,  ��  bx  ��  c@  ��  c@  ��  bx  ��  bx      H   ,  �,  ^�  �,  _X  ��  _X  ��  ^�  �,  ^�      H   ,  ��  `�  ��  a�  ��  a�  ��  `�  ��  `�      H   ,  ��  ^�  ��  _X  ��  _X  ��  ^�  ��  ^�      H   ,  ��  ]   ��  ]�  ��  ]�  ��  ]   ��  ]       H   ,  ��  `   ��  `�  ��  `�  ��  `   ��  `       H   ,  �d  a�  �d  bx  �,  bx  �,  a�  �d  a�      H   ,  ��  ]�  ��  ^�  ��  ^�  ��  ]�  ��  ]�      H   ,  ��  _X  ��  `   ��  `   ��  _X  ��  _X      H   ,  �,  `�  �,  a�  ��  a�  ��  `�  �,  `�      H   ,  ��  ^�  ��  _X  ��  _X  ��  ^�  ��  ^�      H   ,  ��  ]�  ��  ^�  ��  ^�  ��  ]�  ��  ]�      H   ,  ��  ]   ��  ]�  ��  ]�  ��  ]   ��  ]       H   ,  �,  ]�  �,  ^�  ��  ^�  ��  ]�  �,  ]�      H   ,  �d  bx  �d  c@  �,  c@  �,  bx  �d  bx      H   ,  ��  bx  ��  c@  ��  c@  ��  bx  ��  bx      H   ,  ��  a�  ��  bx  �L  bx  �L  a�  ��  a�      H   ,  �,  ]   �,  ]�  ��  ]�  ��  ]   �,  ]       H   ,  ��  ^�  ��  _X  ��  _X  ��  ^�  ��  ^�      H   ,  �,  ]   �,  ]�  ��  ]�  ��  ]   �,  ]       H   ,  ��  `�  ��  a�  ��  a�  ��  `�  ��  `�      H   ,  ��  ]�  ��  ^�  ��  ^�  ��  ]�  ��  ]�      H   ,  ��  _X  ��  `   ��  `   ��  _X  ��  _X      H   ,  ��  ]   ��  ]�  ��  ]�  ��  ]   ��  ]       H   ,  ��  `   ��  `�  ��  `�  ��  `   ��  `       H   ,  ��  N�  ��  O�  �|  O�  �|  N�  ��  N�      H   ,  �l  N�  �l  O�  �4  O�  �4  N�  �l  N�      H   ,  ��  N�  ��  O�  �d  O�  �d  N�  ��  N�      H   ,  �T  N�  �T  O�  �  O�  �  N�  �T  N�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �  N�  �  O�  ��  O�  ��  N�  �  N�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �  N�  �  O�  ��  O�  ��  N�  �  N�      H   ,  ��  S�  ��  Th  �t  Th  �t  S�  ��  S�      H   ,  ��  R�  ��  S�  �t  S�  �t  R�  ��  R�      H   ,  ��  R  ��  R�  �t  R�  �t  R  ��  R      H   ,  ��  QH  ��  R  �t  R  �t  QH  ��  QH      H   ,  ��  P�  ��  QH  �t  QH  �t  P�  ��  P�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  ��  O�  ��  P�  �t  P�  �t  O�  ��  O�      H   ,  ��  L�  ��  M`  �t  M`  �t  L�  ��  L�      H   ,  ��  K�  ��  L�  �t  L�  �t  K�  ��  K�      H   ,  ��  K  ��  K�  �t  K�  �t  K  ��  K      H   ,  ��  J@  ��  K  �t  K  �t  J@  ��  J@      H   ,  ��  Ix  ��  J@  �t  J@  �t  Ix  ��  Ix      H   ,  ��  H�  ��  Ix  �t  Ix  �t  H�  ��  H�      H   ,  �|  N�  �|  O�  �D  O�  �D  N�  �|  N�      H   ,  �  N�  �  O�  ��  O�  ��  N�  �  N�      H   ,  ��  G�  ��  H�  �t  H�  �t  G�  ��  G�      H   ,  ��  G   ��  G�  �t  G�  �t  G   ��  G       H   ,  �d  N�  �d  O�  �,  O�  �,  N�  �d  N�      H   ,  ��  FX  ��  G   �t  G   �t  FX  ��  FX      H   ,  ��  E�  ��  FX  �t  FX  �t  E�  ��  E�      H   ,  ��  D�  ��  E�  �t  E�  �t  D�  ��  D�      H   ,  ��  D   ��  D�  �t  D�  �t  D   ��  D       H   ,  ��  N�  ��  O�  �\  O�  �\  N�  ��  N�      H   ,  ��  C8  ��  D   �t  D   �t  C8  ��  C8      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �$  N�  �$  O�  ��  O�  ��  N�  �$  N�      H   ,  �4  N�  �4  O�  ��  O�  ��  N�  �4  N�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �\  N�  �\  O�  �$  O�  �$  N�  �\  N�      H   ,  �D  N�  �D  O�  �  O�  �  N�  �D  N�      H   ,  ��  N�  ��  O�  �T  O�  �T  N�  ��  N�      H   ,  �,  N�  �,  O�  ��  O�  ��  N�  �,  N�      H   ,  ��  U�  ��  V�  �d  V�  �d  U�  ��  U�      H   ,  ��  P�  ��  QH  �|  QH  �|  P�  ��  P�      H   ,  ��  O�  ��  P�  �|  P�  �|  O�  ��  O�      H   ,  �d  U�  �d  V�  �,  V�  �,  U�  �d  U�      H   ,  ��  R�  ��  S�  �|  S�  �|  R�  ��  R�      H   ,  ��  R  ��  R�  �|  R�  �|  R  ��  R      H   ,  ��  U�  ��  V�  ��  V�  ��  U�  ��  U�      H   ,  �,  U�  �,  V�  ��  V�  ��  U�  �,  U�      H   ,  ��  QH  ��  R  �|  R  �|  QH  ��  QH      H   ,  �d  W�  �d  XP  �,  XP  �,  W�  �d  W�      H   ,  �d  V�  �d  W�  �,  W�  �,  V�  �d  V�      H   ,  ��  Z�  ��  [p  ��  [p  ��  Z�  ��  Z�      H   ,  �d  Y�  �d  Z�  �,  Z�  �,  Y�  �d  Y�      H   ,  ��  W�  ��  XP  �d  XP  �d  W�  ��  W�      H   ,  ��  Y  ��  Y�  ��  Y�  ��  Y  ��  Y      H   ,  ��  XP  ��  Y  ��  Y  ��  XP  ��  XP      H   ,  ��  W�  ��  XP  ��  XP  ��  W�  ��  W�      H   ,  ��  Y�  ��  Z�  ��  Z�  ��  Y�  ��  Y�      H   ,  ��  V�  ��  W�  ��  W�  ��  V�  ��  V�      H   ,  �d  Y  �d  Y�  �,  Y�  �,  Y  �d  Y      H   ,  ��  V�  ��  W�  �d  W�  �d  V�  ��  V�      H   ,  �,  \8  �,  ]   ��  ]   ��  \8  �,  \8      H   ,  �,  [p  �,  \8  ��  \8  ��  [p  �,  [p      H   ,  �,  Z�  �,  [p  ��  [p  ��  Z�  �,  Z�      H   ,  �,  Y�  �,  Z�  ��  Z�  ��  Y�  �,  Y�      H   ,  �,  Y  �,  Y�  ��  Y�  ��  Y  �,  Y      H   ,  ��  \8  ��  ]   ��  ]   ��  \8  ��  \8      H   ,  �,  XP  �,  Y  ��  Y  ��  XP  �,  XP      H   ,  �,  W�  �,  XP  ��  XP  ��  W�  �,  W�      H   ,  �,  V�  �,  W�  ��  W�  ��  V�  �,  V�      H   ,  �d  Z�  �d  [p  �,  [p  �,  Z�  �d  Z�      H   ,  ��  [p  ��  \8  ��  \8  ��  [p  ��  [p      H   ,  �d  XP  �d  Y  �,  Y  �,  XP  �d  XP      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  P�  ��  QH  �\  QH  �\  P�  ��  P�      H   ,  �$  P�  �$  QH  ��  QH  ��  P�  �$  P�      H   ,  �$  QH  �$  R  ��  R  ��  QH  �$  QH      H   ,  ��  O�  ��  P�  �\  P�  �\  O�  ��  O�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  �$  R  �$  R�  ��  R�  ��  R  �$  R      H   ,  �  R�  �  S�  ��  S�  ��  R�  �  R�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �  R  �  R�  ��  R�  ��  R  �  R      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  �$  O�  �$  P�  ��  P�  ��  O�  �$  O�      H   ,  �  QH  �  R  ��  R  ��  QH  �  QH      H   ,  �<  QH  �<  R  �  R  �  QH  �<  QH      H   ,  �<  S�  �<  Th  �  Th  �  S�  �<  S�      H   ,  �<  P�  �<  QH  �  QH  �  P�  �<  P�      H   ,  �$  R�  �$  S�  ��  S�  ��  R�  �$  R�      H   ,  �  P�  �  QH  ��  QH  ��  P�  �  P�      H   ,  �t  S�  �t  Th  �<  Th  �<  S�  �t  S�      H   ,  �  O�  �  P�  ��  P�  ��  O�  �  O�      H   ,  �t  R�  �t  S�  �<  S�  �<  R�  �t  R�      H   ,  ��  S�  ��  Th  �\  Th  �\  S�  ��  S�      H   ,  �t  R  �t  R�  �<  R�  �<  R  �t  R      H   ,  �<  O�  �<  P�  �  P�  �  O�  �<  O�      H   ,  �t  QH  �t  R  �<  R  �<  QH  �t  QH      H   ,  �<  R�  �<  S�  �  S�  �  R�  �<  R�      H   ,  �  S�  �  Th  ��  Th  ��  S�  �  S�      H   ,  ��  R�  ��  S�  �\  S�  �\  R�  ��  R�      H   ,  �t  P�  �t  QH  �<  QH  �<  P�  �t  P�      H   ,  �\  S�  �\  Th  �$  Th  �$  S�  �\  S�      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  �t  O�  �t  P�  �<  P�  �<  O�  �t  O�      H   ,  �\  R�  �\  S�  �$  S�  �$  R�  �\  R�      H   ,  ��  R  ��  R�  �\  R�  �\  R  ��  R      H   ,  �\  R  �\  R�  �$  R�  �$  R  �\  R      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �\  QH  �\  R  �$  R  �$  QH  �\  QH      H   ,  �\  P�  �\  QH  �$  QH  �$  P�  �\  P�      H   ,  �\  O�  �\  P�  �$  P�  �$  O�  �\  O�      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  QH  ��  R  �\  R  �\  QH  ��  QH      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  �<  R  �<  R�  �  R�  �  R  �<  R      H   ,  �d  R  �d  R�  �,  R�  �,  R  �d  R      H   ,  ��  Th  ��  U0  ��  U0  ��  Th  ��  Th      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �  QH  �  R  ��  R  ��  QH  �  QH      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  �  P�  �  QH  ��  QH  ��  P�  �  P�      H   ,  �|  O�  �|  P�  �D  P�  �D  O�  �|  O�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �d  QH  �d  R  �,  R  �,  QH  �d  QH      H   ,  ��  P�  ��  QH  �d  QH  �d  P�  ��  P�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ��  O�  ��  P�  �d  P�  �d  O�  ��  O�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  �d  P�  �d  QH  �,  QH  �,  P�  �d  P�      H   ,  ��  U0  ��  U�  �d  U�  �d  U0  ��  U0      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  ��  U0  ��  U�  ��  U�  ��  U0  ��  U0      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  �d  O�  �d  P�  �,  P�  �,  O�  �d  O�      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  S�  ��  Th  �d  Th  �d  S�  ��  S�      H   ,  ��  R�  ��  S�  �d  S�  �d  R�  ��  R�      H   ,  �  O�  �  P�  ��  P�  ��  O�  �  O�      H   ,  ��  Th  ��  U0  ��  U0  ��  Th  ��  Th      H   ,  �d  U0  �d  U�  �,  U�  �,  U0  �d  U0      H   ,  ��  R  ��  R�  �d  R�  �d  R  ��  R      H   ,  �  R�  �  S�  ��  S�  ��  R�  �  R�      H   ,  �|  R�  �|  S�  �D  S�  �D  R�  �|  R�      H   ,  �d  Th  �d  U0  �,  U0  �,  Th  �d  Th      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  Th  ��  U0  �d  U0  �d  Th  ��  Th      H   ,  �|  R  �|  R�  �D  R�  �D  R  �|  R      H   ,  �d  S�  �d  Th  �,  Th  �,  S�  �d  S�      H   ,  �,  U0  �,  U�  ��  U�  ��  U0  �,  U0      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  �D  R�  �D  S�  �  S�  �  R�  �D  R�      H   ,  �,  Th  �,  U0  ��  U0  ��  Th  �,  Th      H   ,  �|  QH  �|  R  �D  R  �D  QH  �|  QH      H   ,  �D  R  �D  R�  �  R�  �  R  �D  R      H   ,  �,  S�  �,  Th  ��  Th  ��  S�  �,  S�      H   ,  �d  R�  �d  S�  �,  S�  �,  R�  �d  R�      H   ,  �D  QH  �D  R  �  R  �  QH  �D  QH      H   ,  �,  R�  �,  S�  ��  S�  ��  R�  �,  R�      H   ,  �D  P�  �D  QH  �  QH  �  P�  �D  P�      H   ,  �,  R  �,  R�  ��  R�  ��  R  �,  R      H   ,  �D  O�  �D  P�  �  P�  �  O�  �D  O�      H   ,  �,  QH  �,  R  ��  R  ��  QH  �,  QH      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �,  P�  �,  QH  ��  QH  ��  P�  �,  P�      H   ,  �,  O�  �,  P�  ��  P�  ��  O�  �,  O�      H   ,  ��  QH  ��  R  �d  R  �d  QH  ��  QH      H   ,  �|  P�  �|  QH  �D  QH  �D  P�  �|  P�      H   ,  ��  U0  ��  U�  ��  U�  ��  U0  ��  U0      H   ,  �  R  �  R�  ��  R�  ��  R  �  R      H   ,  �  U�  �  V�  ��  V�  ��  U�  �  U�      H   ,  ��  U�  ��  V�  �l  V�  �l  U�  ��  U�      H   ,  ��  R  ��  R�  �l  R�  �l  R  ��  R      H   ,  ��  QH  ��  R  �l  R  �l  QH  ��  QH      H   ,  ��  U0  ��  U�  �l  U�  �l  U0  ��  U0      H   ,  ��  W�  ��  XP  �l  XP  �l  W�  ��  W�      H   ,  ��  P�  ��  QH  �l  QH  �l  P�  ��  P�      H   ,  ��  U�  ��  V�  ��  V�  ��  U�  ��  U�      H   ,  ��  Th  ��  U0  �l  U0  �l  Th  ��  Th      H   ,  �L  U�  �L  V�  �  V�  �  U�  �L  U�      H   ,  ��  R�  ��  S�  �l  S�  �l  R�  ��  R�      H   ,  ��  V�  ��  W�  �l  W�  �l  V�  ��  V�      H   ,  ��  O�  ��  P�  �l  P�  �l  O�  ��  O�      H   ,  ��  U�  ��  V�  �L  V�  �L  U�  ��  U�      H   ,  ��  S�  ��  Th  �l  Th  �l  S�  ��  S�      H   ,  ��  U�  ��  V�  ��  V�  ��  U�  ��  U�      H   ,  �l  U�  �l  V�  �4  V�  �4  U�  �l  U�      H   ,  �l  V�  �l  W�  �4  W�  �4  V�  �l  V�      H   ,  ��  Y  ��  Y�  �L  Y�  �L  Y  ��  Y      H   ,  ��  Y  ��  Y�  ��  Y�  ��  Y  ��  Y      H   ,  �L  Z�  �L  [p  �  [p  �  Z�  �L  Z�      H   ,  ��  XP  ��  Y  ��  Y  ��  XP  ��  XP      H   ,  ��  W�  ��  XP  ��  XP  ��  W�  ��  W�      H   ,  �L  Y�  �L  Z�  �  Z�  �  Y�  �L  Y�      H   ,  ��  V�  ��  W�  ��  W�  ��  V�  ��  V�      H   ,  ��  V�  ��  W�  ��  W�  ��  V�  ��  V�      H   ,  ��  XP  ��  Y  ��  Y  ��  XP  ��  XP      H   ,  ��  \8  ��  ]   ��  ]   ��  \8  ��  \8      H   ,  ��  [p  ��  \8  ��  \8  ��  [p  ��  [p      H   ,  ��  Z�  ��  [p  ��  [p  ��  Z�  ��  Z�      H   ,  �  Y�  �  Z�  ��  Z�  ��  Y�  �  Y�      H   ,  �L  Y  �L  Y�  �  Y�  �  Y  �L  Y      H   ,  ��  Y�  ��  Z�  ��  Z�  ��  Y�  ��  Y�      H   ,  ��  Y  ��  Y�  ��  Y�  ��  Y  ��  Y      H   ,  �L  XP  �L  Y  �  Y  �  XP  �L  XP      H   ,  ��  XP  ��  Y  ��  Y  ��  XP  ��  XP      H   ,  ��  W�  ��  XP  ��  XP  ��  W�  ��  W�      H   ,  �L  W�  �L  XP  �  XP  �  W�  �L  W�      H   ,  ��  V�  ��  W�  ��  W�  ��  V�  ��  V�      H   ,  �L  V�  �L  W�  �  W�  �  V�  �L  V�      H   ,  ��  V�  ��  W�  �L  W�  �L  V�  ��  V�      H   ,  ��  Z�  ��  [p  ��  [p  ��  Z�  ��  Z�      H   ,  ��  [p  ��  \8  ��  \8  ��  [p  ��  [p      H   ,  �  Y  �  Y�  ��  Y�  ��  Y  �  Y      H   ,  �  XP  �  Y  ��  Y  ��  XP  �  XP      H   ,  ��  Y�  ��  Z�  ��  Z�  ��  Y�  ��  Y�      H   ,  �d  \8  �d  ]   �,  ]   �,  \8  �d  \8      H   ,  ��  W�  ��  XP  �L  XP  �L  W�  ��  W�      H   ,  �,  \8  �,  ]   ��  ]   ��  \8  �,  \8      H   ,  �d  [p  �d  \8  �,  \8  �,  [p  �d  [p      H   ,  ��  XP  ��  Y  �L  Y  �L  XP  ��  XP      H   ,  �d  Z�  �d  [p  �,  [p  �,  Z�  �d  Z�      H   ,  �,  [p  �,  \8  ��  \8  ��  [p  �,  [p      H   ,  �d  Y�  �d  Z�  �,  Z�  �,  Y�  �d  Y�      H   ,  �,  Z�  �,  [p  ��  [p  ��  Z�  �,  Z�      H   ,  ��  W�  ��  XP  ��  XP  ��  W�  ��  W�      H   ,  �d  Y  �d  Y�  �,  Y�  �,  Y  �d  Y      H   ,  ��  Y  ��  Y�  ��  Y�  ��  Y  ��  Y      H   ,  �,  Y�  �,  Z�  ��  Z�  ��  Y�  �,  Y�      H   ,  ��  Y�  ��  Z�  �L  Z�  �L  Y�  ��  Y�      H   ,  ��  \8  ��  ]   ��  ]   ��  \8  ��  \8      H   ,  �,  Y  �,  Y�  ��  Y�  ��  Y  �,  Y      H   ,  �,  XP  �,  Y  ��  Y  ��  XP  �,  XP      H   ,  �  W�  �  XP  ��  XP  ��  W�  �  W�      H   ,  ��  \8  ��  ]   �L  ]   �L  \8  ��  \8      H   ,  ��  [p  ��  \8  �L  \8  �L  [p  ��  [p      H   ,  �  V�  �  W�  ��  W�  ��  V�  �  V�      H   ,  ��  Z�  ��  [p  �L  [p  �L  Z�  ��  Z�      H   ,  �L  [p  �L  \8  �  \8  �  [p  �L  [p      H   ,  ��  R�  ��  S�  �L  S�  �L  R�  ��  R�      H   ,  �,  P�  �,  QH  ��  QH  ��  P�  �,  P�      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  �L  U0  �L  U�  �  U�  �  U0  �L  U0      H   ,  �  O�  �  P�  ��  P�  ��  O�  �  O�      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  ��  Th  ��  U0  �L  U0  �L  Th  ��  Th      H   ,  ��  R  ��  R�  �L  R�  �L  R  ��  R      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  �L  Th  �L  U0  �  U0  �  Th  �L  Th      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �L  S�  �L  Th  �  Th  �  S�  �L  S�      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �  QH  �  R  ��  R  ��  QH  �  QH      H   ,  ��  Th  ��  U0  ��  U0  ��  Th  ��  Th      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  �L  R�  �L  S�  �  S�  �  R�  �L  R�      H   ,  ��  QH  ��  R  �L  R  �L  QH  ��  QH      H   ,  �,  R�  �,  S�  ��  S�  ��  R�  �,  R�      H   ,  ��  U0  ��  U�  ��  U�  ��  U0  ��  U0      H   ,  �L  R  �L  R�  �  R�  �  R  �L  R      H   ,  �,  QH  �,  R  ��  R  ��  QH  �,  QH      H   ,  ��  Th  ��  U0  ��  U0  ��  Th  ��  Th      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �L  QH  �L  R  �  R  �  QH  �L  QH      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �  P�  �  QH  ��  QH  ��  P�  �  P�      H   ,  �  U0  �  U�  ��  U�  ��  U0  �  U0      H   ,  �  Th  �  U0  ��  U0  ��  Th  �  Th      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  P�  ��  QH  �L  QH  �L  P�  ��  P�      H   ,  �L  P�  �L  QH  �  QH  �  P�  �L  P�      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �d  Th  �d  U0  �,  U0  �,  Th  �d  Th      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  �  S�  �  Th  ��  Th  ��  S�  �  S�      H   ,  ��  U0  ��  U�  �L  U�  �L  U0  ��  U0      H   ,  �d  S�  �d  Th  �,  Th  �,  S�  �d  S�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  �d  R�  �d  S�  �,  S�  �,  R�  �d  R�      H   ,  ��  O�  ��  P�  �L  P�  �L  O�  ��  O�      H   ,  �d  R  �d  R�  �,  R�  �,  R  �d  R      H   ,  �,  Th  �,  U0  ��  U0  ��  Th  �,  Th      H   ,  �d  QH  �d  R  �,  R  �,  QH  �d  QH      H   ,  �d  P�  �d  QH  �,  QH  �,  P�  �d  P�      H   ,  �,  S�  �,  Th  ��  Th  ��  S�  �,  S�      H   ,  �  R�  �  S�  ��  S�  ��  R�  �  R�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  �L  O�  �L  P�  �  P�  �  O�  �L  O�      H   ,  �  R  �  R�  ��  R�  ��  R  �  R      H   ,  ��  S�  ��  Th  �L  Th  �L  S�  ��  S�      H   ,  �,  R  �,  R�  ��  R�  ��  R  �,  R      H   ,  ��  Th  ��  U0  ��  U0  ��  Th  ��  Th      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �4  O�  �4  P�  ��  P�  ��  O�  �4  O�      H   ,  �T  S�  �T  Th  �  Th  �  S�  �T  S�      H   ,  �4  R  �4  R�  ��  R�  ��  R  �4  R      H   ,  �  S�  �  Th  ��  Th  ��  S�  �  S�      H   ,  �  R  �  R�  ��  R�  ��  R  �  R      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  �l  S�  �l  Th  �4  Th  �4  S�  �l  S�      H   ,  �l  QH  �l  R  �4  R  �4  QH  �l  QH      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  �  O�  �  P�  ��  P�  ��  O�  �  O�      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  �l  U0  �l  U�  �4  U�  �4  U0  �l  U0      H   ,  �T  P�  �T  QH  �  QH  �  P�  �T  P�      H   ,  �  R�  �  S�  ��  S�  ��  R�  �  R�      H   ,  �4  QH  �4  R  ��  R  ��  QH  �4  QH      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  �4  U0  �4  U�  ��  U�  ��  U0  �4  U0      H   ,  �T  R  �T  R�  �  R�  �  R  �T  R      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �4  Th  �4  U0  ��  U0  ��  Th  �4  Th      H   ,  ��  S�  ��  Th  �T  Th  �T  S�  ��  S�      H   ,  �l  Th  �l  U0  �4  U0  �4  Th  �l  Th      H   ,  �  QH  �  R  ��  R  ��  QH  �  QH      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ��  R�  ��  S�  �T  S�  �T  R�  ��  R�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �l  P�  �l  QH  �4  QH  �4  P�  �l  P�      H   ,  �T  O�  �T  P�  �  P�  �  O�  �T  O�      H   ,  ��  R  ��  R�  �T  R�  �T  R  ��  R      H   ,  �l  R  �l  R�  �4  R�  �4  R  �l  R      H   ,  �4  S�  �4  Th  ��  Th  ��  S�  �4  S�      H   ,  ��  QH  ��  R  �T  R  �T  QH  ��  QH      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  �T  QH  �T  R  �  R  �  QH  �T  QH      H   ,  ��  P�  ��  QH  �T  QH  �T  P�  ��  P�      H   ,  �l  O�  �l  P�  �4  P�  �4  O�  �l  O�      H   ,  �l  R�  �l  S�  �4  S�  �4  R�  �l  R�      H   ,  ��  O�  ��  P�  �T  P�  �T  O�  ��  O�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �4  P�  �4  QH  ��  QH  ��  P�  �4  P�      H   ,  ��  Th  ��  U0  ��  U0  ��  Th  ��  Th      H   ,  �  P�  �  QH  ��  QH  ��  P�  �  P�      H   ,  �4  R�  �4  S�  ��  S�  ��  R�  �4  R�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �T  R�  �T  S�  �  S�  �  R�  �T  R�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  �T  G�  �T  H�  �  H�  �  G�  �T  G�      H   ,  ��  K  ��  K�  ��  K�  ��  K  ��  K      H   ,  ��  H�  ��  Ix  ��  Ix  ��  H�  ��  H�      H   ,  ��  FX  ��  G   ��  G   ��  FX  ��  FX      H   ,  ��  J@  ��  K  ��  K  ��  J@  ��  J@      H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  �T  G   �T  G�  �  G�  �  G   �T  G       H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �  G   �  G�  ��  G�  ��  G   �  G       H   ,  ��  G�  ��  H�  ��  H�  ��  G�  ��  G�      H   ,  �  J@  �  K  ��  K  ��  J@  �  J@      H   ,  �  L�  �  M`  ��  M`  ��  L�  �  L�      H   ,  �  FX  �  G   ��  G   ��  FX  �  FX      H   ,  �4  N(  �4  N�  ��  N�  ��  N(  �4  N(      H   ,  ��  E�  ��  FX  ��  FX  ��  E�  ��  E�      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  ��  Ix  ��  J@  ��  J@  ��  Ix  ��  Ix      H   ,  �4  M`  �4  N(  ��  N(  ��  M`  �4  M`      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  �  Ix  �  J@  ��  J@  ��  Ix  �  Ix      H   ,  �T  K  �T  K�  �  K�  �  K  �T  K      H   ,  �  E�  �  FX  ��  FX  ��  E�  �  E�      H   ,  �4  L�  �4  M`  ��  M`  ��  L�  �4  L�      H   ,  �T  M`  �T  N(  �  N(  �  M`  �T  M`      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �l  N(  �l  N�  �4  N�  �4  N(  �l  N(      H   ,  �  K�  �  L�  ��  L�  ��  K�  �  K�      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  �T  K�  �T  L�  �  L�  �  K�  �T  K�      H   ,  �  N(  �  N�  ��  N�  ��  N(  �  N(      H   ,  �  H�  �  Ix  ��  Ix  ��  H�  �  H�      H   ,  �T  J@  �T  K  �  K  �  J@  �T  J@      H   ,  ��  D�  ��  E�  ��  E�  ��  D�  ��  D�      H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  �T  N(  �T  N�  �  N�  �  N(  �T  N(      H   ,  ��  G   ��  G�  ��  G�  ��  G   ��  G       H   ,  �  K  �  K�  ��  K�  ��  K  �  K      H   ,  ��  J@  ��  K  ��  K  ��  J@  ��  J@      H   ,  �T  Ix  �T  J@  �  J@  �  Ix  �T  Ix      H   ,  ��  N(  ��  N�  �T  N�  �T  N(  ��  N(      H   ,  ��  M`  ��  N(  �T  N(  �T  M`  ��  M`      H   ,  ��  L�  ��  M`  �T  M`  �T  L�  ��  L�      H   ,  ��  K�  ��  L�  �T  L�  �T  K�  ��  K�      H   ,  ��  K  ��  K�  �T  K�  �T  K  ��  K      H   ,  ��  J@  ��  K  �T  K  �T  J@  ��  J@      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  ��  Ix  ��  J@  �T  J@  �T  Ix  ��  Ix      H   ,  ��  K  ��  K�  ��  K�  ��  K  ��  K      H   ,  ��  H�  ��  Ix  �T  Ix  �T  H�  ��  H�      H   ,  �  M`  �  N(  ��  N(  ��  M`  �  M`      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �T  H�  �T  Ix  �  Ix  �  H�  �T  H�      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  �T  L�  �T  M`  �  M`  �  L�  �T  L�      H   ,  �  G�  �  H�  ��  H�  ��  G�  �  G�      H   ,  ��  J@  ��  K  �|  K  �|  J@  ��  J@      H   ,  ��  C8  ��  D   �|  D   �|  C8  ��  C8      H   ,  ��  H�  ��  Ix  �|  Ix  �|  H�  ��  H�      H   ,  ��  G�  ��  H�  ��  H�  ��  G�  ��  G�      H   ,  ��  E�  ��  FX  �|  FX  �|  E�  ��  E�      H   ,  ��  Bp  ��  C8  �|  C8  �|  Bp  ��  Bp      H   ,  �$  G�  �$  H�  ��  H�  ��  G�  �$  G�      H   ,  �|  G�  �|  H�  �D  H�  �D  G�  �|  G�      H   ,  ��  G�  ��  H�  ��  H�  ��  G�  ��  G�      H   ,  ��  Ix  ��  J@  �|  J@  �|  Ix  ��  Ix      H   ,  ��  A�  ��  Bp  �|  Bp  �|  A�  ��  A�      H   ,  ��  G   ��  G�  �|  G�  �|  G   ��  G       H   ,  ��  D�  ��  E�  �|  E�  �|  D�  ��  D�      H   ,  �  G�  �  H�  ��  H�  ��  G�  �  G�      H   ,  �<  G�  �<  H�  �  H�  �  G�  �<  G�      H   ,  ��  K  ��  K�  �|  K�  �|  K  ��  K      H   ,  �t  G�  �t  H�  �<  H�  �<  G�  �t  G�      H   ,  ��  K�  ��  L�  �|  L�  �|  K�  ��  K�      H   ,  ��  FX  ��  G   �|  G   �|  FX  ��  FX      H   ,  ��  D   ��  D�  �|  D�  �|  D   ��  D       H   ,  �  G�  �  H�  ��  H�  ��  G�  �  G�      H   ,  �D  G�  �D  H�  �  H�  �  G�  �D  G�      H   ,  ��  G�  ��  H�  �|  H�  �|  G�  ��  G�      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  ��  Ix  ��  J@  �d  J@  �d  Ix  ��  Ix      H   ,  �d  M`  �d  N(  �,  N(  �,  M`  �d  M`      H   ,  �  J@  �  K  ��  K  ��  J@  �  J@      H   ,  �|  J@  �|  K  �D  K  �D  J@  �|  J@      H   ,  �d  K�  �d  L�  �,  L�  �,  K�  �d  K�      H   ,  �  Ix  �  J@  ��  J@  ��  Ix  �  Ix      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  ��  N(  ��  N�  �d  N�  �d  N(  ��  N(      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  �  H�  �  Ix  ��  Ix  ��  H�  �  H�      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  ��  H�  ��  Ix  ��  Ix  ��  H�  ��  H�      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  ��  K�  ��  L�  �d  L�  �d  K�  ��  K�      H   ,  ��  L�  ��  M`  �d  M`  �d  L�  ��  L�      H   ,  �|  Ix  �|  J@  �D  J@  �D  Ix  �|  Ix      H   ,  �  K  �  K�  ��  K�  ��  K  �  K      H   ,  �|  K�  �|  L�  �D  L�  �D  K�  �|  K�      H   ,  ��  K  ��  K�  ��  K�  ��  K  ��  K      H   ,  �  M`  �  N(  ��  N(  ��  M`  �  M`      H   ,  �|  N(  �|  N�  �D  N�  �D  N(  �|  N(      H   ,  �|  H�  �|  Ix  �D  Ix  �D  H�  �|  H�      H   ,  �D  N(  �D  N�  �  N�  �  N(  �D  N(      H   ,  �|  K  �|  K�  �D  K�  �D  K  �|  K      H   ,  �  L�  �  M`  ��  M`  ��  L�  �  L�      H   ,  �D  M`  �D  N(  �  N(  �  M`  �D  M`      H   ,  �D  L�  �D  M`  �  M`  �  L�  �D  L�      H   ,  �,  N(  �,  N�  ��  N�  ��  N(  �,  N(      H   ,  ��  J@  ��  K  ��  K  ��  J@  ��  J@      H   ,  �D  K�  �D  L�  �  L�  �  K�  �D  K�      H   ,  �,  M`  �,  N(  ��  N(  ��  M`  �,  M`      H   ,  �D  K  �D  K�  �  K�  �  K  �D  K      H   ,  �D  J@  �D  K  �  K  �  J@  �D  J@      H   ,  �|  M`  �|  N(  �D  N(  �D  M`  �|  M`      H   ,  �D  Ix  �D  J@  �  J@  �  Ix  �D  Ix      H   ,  ��  K  ��  K�  �d  K�  �d  K  ��  K      H   ,  �D  H�  �D  Ix  �  Ix  �  H�  �D  H�      H   ,  �  K�  �  L�  ��  L�  ��  K�  �  K�      H   ,  ��  M`  ��  N(  �d  N(  �d  M`  ��  M`      H   ,  �d  L�  �d  M`  �,  M`  �,  L�  �d  L�      H   ,  ��  J@  ��  K  �d  K  �d  J@  ��  J@      H   ,  �|  L�  �|  M`  �D  M`  �D  L�  �|  L�      H   ,  �d  N(  �d  N�  �,  N�  �,  N(  �d  N(      H   ,  ��  Ix  ��  J@  ��  J@  ��  Ix  ��  Ix      H   ,  �  N(  �  N�  ��  N�  ��  N(  �  N(      H   ,  �t  Ix  �t  J@  �<  J@  �<  Ix  �t  Ix      H   ,  �t  K  �t  K�  �<  K�  �<  K  �t  K      H   ,  �<  H�  �<  Ix  �  Ix  �  H�  �<  H�      H   ,  ��  Ix  ��  J@  ��  J@  ��  Ix  ��  Ix      H   ,  �t  J@  �t  K  �<  K  �<  J@  �t  J@      H   ,  �t  H�  �t  Ix  �<  Ix  �<  H�  �t  H�      H   ,  ��  H�  ��  Ix  ��  Ix  ��  H�  ��  H�      H   ,  �<  Ix  �<  J@  �  J@  �  Ix  �<  Ix      H   ,  �  FX  �  G   ��  G   ��  FX  �  FX      H   ,  �$  A�  �$  Bp  ��  Bp  ��  A�  �$  A�      H   ,  ��  Bp  ��  C8  ��  C8  ��  Bp  ��  Bp      H   ,  �<  A�  �<  Bp  �  Bp  �  A�  �<  A�      H   ,  ��  C8  ��  D   ��  D   ��  C8  ��  C8      H   ,  �<  D   �<  D�  �  D�  �  D   �<  D       H   ,  �t  G   �t  G�  �<  G�  �<  G   �t  G       H   ,  �\  E�  �\  FX  �$  FX  �$  E�  �\  E�      H   ,  ��  E�  ��  FX  ��  FX  ��  E�  ��  E�      H   ,  �  Bp  �  C8  ��  C8  ��  Bp  �  Bp      H   ,  ��  C8  ��  D   ��  D   ��  C8  ��  C8      H   ,  �t  FX  �t  G   �<  G   �<  FX  �t  FX      H   ,  �\  D�  �\  E�  �$  E�  �$  D�  �\  D�      H   ,  �<  FX  �<  G   �  G   �  FX  �<  FX      H   ,  �$  D   �$  D�  ��  D�  ��  D   �$  D       H   ,  �t  E�  �t  FX  �<  FX  �<  E�  �t  E�      H   ,  �\  D   �\  D�  �$  D�  �$  D   �\  D       H   ,  ��  Bp  ��  C8  ��  C8  ��  Bp  ��  Bp      H   ,  �$  G   �$  G�  ��  G�  ��  G   �$  G       H   ,  ��  D�  ��  E�  �\  E�  �\  D�  ��  D�      H   ,  �t  D�  �t  E�  �<  E�  �<  D�  �t  D�      H   ,  �\  C8  �\  D   �$  D   �$  C8  �\  C8      H   ,  ��  C8  ��  D   �\  D   �\  C8  ��  C8      H   ,  �  E�  �  FX  ��  FX  ��  E�  �  E�      H   ,  ��  E�  ��  FX  ��  FX  ��  E�  ��  E�      H   ,  �t  D   �t  D�  �<  D�  �<  D   �t  D       H   ,  �\  Bp  �\  C8  �$  C8  �$  Bp  �\  Bp      H   ,  �  A�  �  Bp  ��  Bp  ��  A�  �  A�      H   ,  ��  A�  ��  Bp  ��  Bp  ��  A�  ��  A�      H   ,  �t  C8  �t  D   �<  D   �<  C8  �t  C8      H   ,  �\  A�  �\  Bp  �$  Bp  �$  A�  �\  A�      H   ,  �<  G   �<  G�  �  G�  �  G   �<  G       H   ,  �  D�  �  E�  ��  E�  ��  D�  �  D�      H   ,  �<  C8  �<  D   �  D   �  C8  �<  C8      H   ,  �t  Bp  �t  C8  �<  C8  �<  Bp  �t  Bp      H   ,  �$  C8  �$  D   ��  D   ��  C8  �$  C8      H   ,  �<  E�  �<  FX  �  FX  �  E�  �<  E�      H   ,  ��  D�  ��  E�  ��  E�  ��  D�  ��  D�      H   ,  �t  A�  �t  Bp  �<  Bp  �<  A�  �t  A�      H   ,  ��  Bp  ��  C8  �\  C8  �\  Bp  ��  Bp      H   ,  ��  FX  ��  G   ��  G   ��  FX  ��  FX      H   ,  ��  A�  ��  Bp  ��  Bp  ��  A�  ��  A�      H   ,  �  D   �  D�  ��  D�  ��  D   �  D       H   ,  ��  D�  ��  E�  ��  E�  ��  D�  ��  D�      H   ,  �<  D�  �<  E�  �  E�  �  D�  �<  D�      H   ,  ��  D   ��  D�  �\  D�  �\  D   ��  D       H   ,  ��  A�  ��  Bp  �\  Bp  �\  A�  ��  A�      H   ,  �<  Bp  �<  C8  �  C8  �  Bp  �<  Bp      H   ,  ��  D   ��  D�  ��  D�  ��  D   ��  D       H   ,  �  G   �  G�  ��  G�  ��  G   �  G       H   ,  �$  E�  �$  FX  ��  FX  ��  E�  �$  E�      H   ,  �$  Bp  �$  C8  ��  C8  ��  Bp  �$  Bp      H   ,  �$  FX  �$  G   ��  G   ��  FX  �$  FX      H   ,  ��  FX  ��  G   ��  G   ��  FX  ��  FX      H   ,  �  C8  �  D   ��  D   ��  C8  �  C8      H   ,  ��  D   ��  D�  ��  D�  ��  D   ��  D       H   ,  �$  D�  �$  E�  ��  E�  ��  D�  �$  D�      H   ,  ��  G   ��  G�  ��  G�  ��  G   ��  G       H   ,  �|  D�  �|  E�  �D  E�  �D  D�  �|  D�      H   ,  �|  A�  �|  Bp  �D  Bp  �D  A�  �|  A�      H   ,  �D  D   �D  D�  �  D�  �  D   �D  D       H   ,  �|  E�  �|  FX  �D  FX  �D  E�  �|  E�      H   ,  �  FX  �  G   ��  G   ��  FX  �  FX      H   ,  �|  Bp  �|  C8  �D  C8  �D  Bp  �|  Bp      H   ,  �D  G   �D  G�  �  G�  �  G   �D  G       H   ,  �  G   �  G�  ��  G�  ��  G   �  G       H   ,  �|  FX  �|  G   �D  G   �D  FX  �|  FX      H   ,  �D  FX  �D  G   �  G   �  FX  �D  FX      H   ,  �|  C8  �|  D   �D  D   �D  C8  �|  C8      H   ,  �  E�  �  FX  ��  FX  ��  E�  �  E�      H   ,  �D  E�  �D  FX  �  FX  �  E�  �D  E�      H   ,  ��  G   ��  G�  ��  G�  ��  G   ��  G       H   ,  �|  D   �|  D�  �D  D�  �D  D   �|  D       H   ,  �D  D�  �D  E�  �  E�  �  D�  �D  D�      H   ,  �|  G   �|  G�  �D  G�  �D  G   �|  G       H   ,  �  K  �  K�  ��  K�  ��  K  �  K      H   ,  �  J@  �  K  ��  K  ��  J@  �  J@      H   ,  �L  N�  �L  O�  �  O�  �  N�  �L  N�      H   ,  �  Ix  �  J@  ��  J@  ��  Ix  �  Ix      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �  H�  �  Ix  ��  Ix  ��  H�  �  H�      H   ,  �  G�  �  H�  ��  H�  ��  G�  �  G�      H   ,  �  G   �  G�  ��  G�  ��  G   �  G       H   ,  �  FX  �  G   ��  G   ��  FX  �  FX      H   ,  ��  N�  ��  O�  �l  O�  �l  N�  ��  N�      H   ,  �  E�  �  FX  ��  FX  ��  E�  �  E�      H   ,  ��  N�  ��  O�  �T  O�  �T  N�  ��  N�      H   ,  �  D�  �  E�  ��  E�  ��  D�  �  D�      H   ,  �4  N�  �4  O�  ��  O�  ��  N�  �4  N�      H   ,  �  D   �  D�  ��  D�  ��  D   �  D       H   ,  �  C8  �  D   ��  D   ��  C8  �  C8      H   ,  ��  N�  ��  O�  ƴ  O�  ƴ  N�  ��  N�      H   ,  �\  N�  �\  O�  �$  O�  �$  N�  �\  N�      H   ,  �  Bp  �  C8  ��  C8  ��  Bp  �  Bp      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �  A�  �  Bp  ��  Bp  ��  A�  �  A�      H   ,  �D  N�  �D  O�  �  O�  �  N�  �D  N�      H   ,  �l  N�  �l  O�  �4  O�  �4  N�  �l  N�      H   ,  �  N�  �  O�  ��  O�  ��  N�  �  N�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  ��  N�  ��  O�  �L  O�  �L  N�  ��  N�      H   ,  �  P�  �  QH  ��  QH  ��  P�  �  P�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  Ô  N�  Ô  O�  �\  O�  �\  N�  Ô  N�      H   ,  �  O�  �  P�  ��  P�  ��  O�  �  O�      H   ,  ƴ  N�  ƴ  O�  �|  O�  �|  N�  ƴ  N�      H   ,  �T  N�  �T  O�  �  O�  �  N�  �T  N�      H   ,  ��  N�  ��  O�  �t  O�  �t  N�  ��  N�      H   ,  �  N�  �  O�  ��  O�  ��  N�  �  N�      H   ,  �<  N�  �<  O�  �  O�  �  N�  �<  N�      H   ,  �$  N�  �$  O�  ��  O�  ��  N�  �$  N�      H   ,  �  N(  �  N�  ��  N�  ��  N(  �  N(      H   ,  ��  N�  ��  O�  Ô  O�  Ô  N�  ��  N�      H   ,  �  M`  �  N(  ��  N(  ��  M`  �  M`      H   ,  �  L�  �  M`  ��  M`  ��  L�  �  L�      H   ,  �  N�  �  O�  ��  O�  ��  N�  �  N�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �t  N�  �t  O�  �<  O�  �<  N�  �t  N�      H   ,  �  K�  �  L�  ��  L�  ��  K�  �  K�      H   ,  �|  N�  �|  O�  �D  O�  �D  N�  �|  N�      H   ,  �$  O�  �$  P�  ��  P�  ��  O�  �$  O�      H   ,  ƴ  O�  ƴ  P�  �|  P�  �|  O�  ƴ  O�      H   ,  ��  P�  ��  QH  ƴ  QH  ƴ  P�  ��  P�      H   ,  ��  O�  ��  P�  Ô  P�  Ô  O�  ��  O�      H   ,  Ô  P�  Ô  QH  �\  QH  �\  P�  Ô  P�      H   ,  �\  O�  �\  P�  �$  P�  �$  O�  �\  O�      H   ,  ��  O�  ��  P�  ƴ  P�  ƴ  O�  ��  O�      H   ,  �\  P�  �\  QH  �$  QH  �$  P�  �\  P�      H   ,  Ô  O�  Ô  P�  �\  P�  �\  O�  Ô  O�      H   ,  ��  P�  ��  QH  Ô  QH  Ô  P�  ��  P�      H   ,  �|  O�  �|  P�  �D  P�  �D  O�  �|  O�      H   ,  �$  P�  �$  QH  ��  QH  ��  P�  �$  P�      H   ,  ƴ  P�  ƴ  QH  �|  QH  �|  P�  ƴ  P�      H   ,  ��  V�  ��  W�  �L  W�  �L  V�  ��  V�      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  ��  U�  ��  V�  �L  V�  �L  U�  ��  U�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  U0  ��  U�  �L  U�  �L  U0  ��  U0      H   ,  �L  [p  �L  \8  �  \8  �  [p  �L  [p      H   ,  ��  R  ��  R�  �L  R�  �L  R  ��  R      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  ��  QH  ��  R  �L  R  �L  QH  ��  QH      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  P�  ��  QH  �L  QH  �L  P�  ��  P�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ��  O�  ��  P�  �L  P�  �L  O�  ��  O�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �<  P�  �<  QH  �  QH  �  P�  �<  P�      H   ,  ��  O�  ��  P�  �l  P�  �l  O�  ��  O�      H   ,  �4  P�  �4  QH  ��  QH  ��  P�  �4  P�      H   ,  ��  O�  ��  P�  �T  P�  �T  O�  ��  O�      H   ,  �L  P�  �L  QH  �  QH  �  P�  �L  P�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  �L  Z�  �L  [p  �  [p  �  Z�  �L  Z�      H   ,  �  \8  �  ]   ��  ]   ��  \8  �  \8      H   ,  �4  O�  �4  P�  ��  P�  ��  O�  �4  O�      H   ,  �  [p  �  \8  ��  \8  ��  [p  �  [p      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �T  O�  �T  P�  �  P�  �  O�  �T  O�      H   ,  ��  O�  ��  P�  �t  P�  �t  O�  ��  O�      H   ,  ��  QH  ��  R  �l  R  �l  QH  ��  QH      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  �L  Y�  �L  Z�  �  Z�  �  Y�  �L  Y�      H   ,  �  Z�  �  [p  ��  [p  ��  Z�  �  Z�      H   ,  ��  \8  ��  ]   ��  ]   ��  \8  ��  \8      H   ,  �<  O�  �<  P�  �  P�  �  O�  �<  O�      H   ,  ��  [p  ��  \8  ��  \8  ��  [p  ��  [p      H   ,  ��  P�  ��  QH  �l  QH  �l  P�  ��  P�      H   ,  �l  P�  �l  QH  �4  QH  �4  P�  �l  P�      H   ,  �  QH  �  R  ��  R  ��  QH  �  QH      H   ,  �l  O�  �l  P�  �4  P�  �4  O�  �l  O�      H   ,  �L  Y  �L  Y�  �  Y�  �  Y  �L  Y      H   ,  ��  \8  ��  ]   �L  ]   �L  \8  ��  \8      H   ,  ��  Z�  ��  [p  ��  [p  ��  Z�  ��  Z�      H   ,  �L  O�  �L  P�  �  P�  �  O�  �L  O�      H   ,  ��  [p  ��  \8  �L  \8  �L  [p  ��  [p      H   ,  ��  Y�  ��  Z�  ��  Z�  ��  Y�  ��  Y�      H   ,  ��  Y  ��  Y�  ��  Y�  ��  Y  ��  Y      H   ,  �  P�  �  QH  ��  QH  ��  P�  �  P�      H   ,  ��  XP  ��  Y  ��  Y  ��  XP  ��  XP      H   ,  �L  XP  �L  Y  �  Y  �  XP  �L  XP      H   ,  ��  Z�  ��  [p  �L  [p  �L  Z�  ��  Z�      H   ,  ��  W�  ��  XP  ��  XP  ��  W�  ��  W�      H   ,  ��  V�  ��  W�  ��  W�  ��  V�  ��  V�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  �L  W�  �L  XP  �  XP  �  W�  �L  W�      H   ,  ��  Y�  ��  Z�  �L  Z�  �L  Y�  ��  Y�      H   ,  ��  U�  ��  V�  ��  V�  ��  U�  ��  U�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  �  O�  �  P�  ��  P�  ��  O�  �  O�      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  U0  ��  U�  ��  U�  ��  U0  ��  U0      H   ,  �L  QH  �L  R  �  R  �  QH  �L  QH      H   ,  �L  \8  �L  ]   �  ]   �  \8  �L  \8      H   ,  �t  O�  �t  P�  �<  P�  �<  O�  �t  O�      H   ,  ��  Y  ��  Y�  �L  Y�  �L  Y  ��  Y      H   ,  �  O�  �  P�  ��  P�  ��  O�  �  O�      H   ,  ��  XP  ��  Y  �L  Y  �L  XP  ��  XP      H   ,  ��  W�  ��  XP  �L  XP  �L  W�  ��  W�      H   ,  ��  Th  ��  U0  ��  U0  ��  Th  ��  Th      H   ,  �<  G�  �<  H�  �  H�  �  G�  �<  G�      H   ,  �  G�  �  H�  ��  H�  ��  G�  �  G�      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  �t  G�  �t  H�  �<  H�  �<  G�  �t  G�      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  �T  G�  �T  H�  �  H�  �  G�  �T  G�      H   ,  ��  G�  ��  H�  �t  H�  �t  G�  ��  G�      H   ,  ��  G�  ��  H�  �T  H�  �T  G�  ��  G�      H   ,  ��  G�  ��  H�  ��  H�  ��  G�  ��  G�      H   ,  ��  K�  ��  L�  �T  L�  �T  K�  ��  K�      H   ,  �<  K  �<  K�  �  K�  �  K  �<  K      H   ,  �t  Ix  �t  J@  �<  J@  �<  Ix  �t  Ix      H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  ��  K  ��  K�  �T  K�  �T  K  ��  K      H   ,  ��  N(  ��  N�  �T  N�  �T  N(  ��  N(      H   ,  ��  M`  ��  N(  �T  N(  �T  M`  ��  M`      H   ,  �t  H�  �t  Ix  �<  Ix  �<  H�  �t  H�      H   ,  ��  N(  ��  N�  �t  N�  �t  N(  ��  N(      H   ,  �T  N(  �T  N�  �  N�  �  N(  �T  N(      H   ,  ��  J@  ��  K  �T  K  �T  J@  ��  J@      H   ,  ��  M`  ��  N(  �t  N(  �t  M`  ��  M`      H   ,  �T  M`  �T  N(  �  N(  �  M`  �T  M`      H   ,  �  J@  �  K  ��  K  ��  J@  �  J@      H   ,  �T  L�  �T  M`  �  M`  �  L�  �T  L�      H   ,  ��  L�  ��  M`  �t  M`  �t  L�  ��  L�      H   ,  �T  K�  �T  L�  �  L�  �  K�  �T  K�      H   ,  ��  K�  ��  L�  �t  L�  �t  K�  ��  K�      H   ,  �T  K  �T  K�  �  K�  �  K  �T  K      H   ,  �<  Ix  �<  J@  �  J@  �  Ix  �<  Ix      H   ,  �T  J@  �T  K  �  K  �  J@  �T  J@      H   ,  ��  K  ��  K�  �t  K�  �t  K  ��  K      H   ,  �T  Ix  �T  J@  �  J@  �  Ix  �T  Ix      H   ,  ��  J@  ��  K  �t  K  �t  J@  ��  J@      H   ,  �T  H�  �T  Ix  �  Ix  �  H�  �T  H�      H   ,  �  Ix  �  J@  ��  J@  ��  Ix  �  Ix      H   ,  ��  L�  ��  M`  �T  M`  �T  L�  ��  L�      H   ,  ��  Ix  ��  J@  �t  J@  �t  Ix  ��  Ix      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  ��  H�  ��  Ix  �t  Ix  �t  H�  ��  H�      H   ,  ��  Ix  ��  J@  �T  J@  �T  Ix  ��  Ix      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �t  J@  �t  K  �<  K  �<  J@  �t  J@      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �<  K�  �<  L�  �  L�  �  K�  �<  K�      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  �<  H�  �<  Ix  �  Ix  �  H�  �<  H�      H   ,  ��  H�  ��  Ix  �T  Ix  �T  H�  ��  H�      H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  ��  K  ��  K�  ��  K�  ��  K  ��  K      H   ,  �  H�  �  Ix  ��  Ix  ��  H�  �  H�      H   ,  �  L�  �  M`  ��  M`  ��  L�  �  L�      H   ,  ��  J@  ��  K  ��  K  ��  J@  ��  J@      H   ,  �  K�  �  L�  ��  L�  ��  K�  �  K�      H   ,  �  K  �  K�  ��  K�  ��  K  �  K      H   ,  �<  J@  �<  K  �  K  �  J@  �<  J@      H   ,  ��  Ix  ��  J@  ��  J@  ��  Ix  ��  Ix      H   ,  �<  N(  �<  N�  �  N�  �  N(  �<  N(      H   ,  ��  H�  ��  Ix  ��  Ix  ��  H�  ��  H�      H   ,  �  N(  �  N�  ��  N�  ��  N(  �  N(      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  �<  M`  �<  N(  �  N(  �  M`  �<  M`      H   ,  �<  L�  �<  M`  �  M`  �  L�  �<  L�      H   ,  �t  N(  �t  N�  �<  N�  �<  N(  �t  N(      H   ,  �t  M`  �t  N(  �<  N(  �<  M`  �t  M`      H   ,  �  M`  �  N(  ��  N(  ��  M`  �  M`      H   ,  �t  L�  �t  M`  �<  M`  �<  L�  �t  L�      H   ,  �t  K  �t  K�  �<  K�  �<  K  �t  K      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  �t  K�  �t  L�  �<  L�  �<  K�  �t  K�      H   ,  �  M`  �  N(  ��  N(  ��  M`  �  M`      H   ,  �4  L�  �4  M`  ��  M`  ��  L�  �4  L�      H   ,  �4  N(  �4  N�  ��  N�  ��  N(  �4  N(      H   ,  �L  N(  �L  N�  �  N�  �  N(  �L  N(      H   ,  ��  N(  ��  N�  �l  N�  �l  N(  ��  N(      H   ,  �4  M`  �4  N(  ��  N(  ��  M`  �4  M`      H   ,  �4  K�  �4  L�  ��  L�  ��  K�  �4  K�      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  ��  N(  ��  N�  �L  N�  �L  N(  ��  N(      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �l  L�  �l  M`  �4  M`  �4  L�  �l  L�      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  ��  M`  ��  N(  �L  N(  �L  M`  ��  M`      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  �l  M`  �l  N(  �4  N(  �4  M`  �l  M`      H   ,  ��  M`  ��  N(  �l  N(  �l  M`  ��  M`      H   ,  ��  L�  ��  M`  �l  M`  �l  L�  ��  L�      H   ,  �l  N(  �l  N�  �4  N�  �4  N(  �l  N(      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �  N(  �  N�  ��  N�  ��  N(  �  N(      H   ,  �L  M`  �L  N(  �  N(  �  M`  �L  M`      H   ,  �t  C8  �t  D   �<  D   �<  C8  �t  C8      H   ,  �T  D�  �T  E�  �  E�  �  D�  �T  D�      H   ,  �t  E�  �t  FX  �<  FX  �<  E�  �t  E�      H   ,  ��  G   ��  G�  �t  G�  �t  G   ��  G       H   ,  �T  D   �T  D�  �  D�  �  D   �T  D       H   ,  ��  G   ��  G�  ��  G�  ��  G   ��  G       H   ,  ��  FX  ��  G   �t  G   �t  FX  ��  FX      H   ,  �<  D   �<  D�  �  D�  �  D   �<  D       H   ,  �<  G   �<  G�  �  G�  �  G   �<  G       H   ,  ��  E�  ��  FX  �t  FX  �t  E�  ��  E�      H   ,  ��  E�  ��  FX  ��  FX  ��  E�  ��  E�      H   ,  �<  Bp  �<  C8  �  C8  �  Bp  �<  Bp      H   ,  ��  D�  ��  E�  �t  E�  �t  D�  ��  D�      H   ,  ��  C8  ��  D   ��  D   ��  C8  ��  C8      H   ,  ��  D   ��  D�  �t  D�  �t  D   ��  D       H   ,  �t  G   �t  G�  �<  G�  �<  G   �t  G       H   ,  �t  D   �t  D�  �<  D�  �<  D   �t  D       H   ,  ��  C8  ��  D   �t  D   �t  C8  ��  C8      H   ,  �t  D�  �t  E�  �<  E�  �<  D�  �t  D�      H   ,  �  D�  �  E�  ��  E�  ��  D�  �  D�      H   ,  ��  Bp  ��  C8  �t  C8  �t  Bp  ��  Bp      H   ,  �<  D�  �<  E�  �  E�  �  D�  �<  D�      H   ,  ��  A�  ��  Bp  �t  Bp  �t  A�  ��  A�      H   ,  �  FX  �  G   ��  G   ��  FX  �  FX      H   ,  �t  A�  �t  Bp  �<  Bp  �<  A�  �t  A�      H   ,  �  G   �  G�  ��  G�  ��  G   �  G       H   ,  ��  E�  ��  FX  �T  FX  �T  E�  ��  E�      H   ,  �<  A�  �<  Bp  �  Bp  �  A�  �<  A�      H   ,  ��  FX  ��  G   �T  G   �T  FX  ��  FX      H   ,  �  C8  �  D   ��  D   ��  C8  �  C8      H   ,  �<  E�  �<  FX  �  FX  �  E�  �<  E�      H   ,  ��  Bp  ��  C8  ��  C8  ��  Bp  ��  Bp      H   ,  ��  D�  ��  E�  ��  E�  ��  D�  ��  D�      H   ,  �  D   �  D�  ��  D�  ��  D   �  D       H   ,  �T  G   �T  G�  �  G�  �  G   �T  G       H   ,  �<  FX  �<  G   �  G   �  FX  �<  FX      H   ,  �t  Bp  �t  C8  �<  C8  �<  Bp  �t  Bp      H   ,  �T  FX  �T  G   �  G   �  FX  �T  FX      H   ,  ��  FX  ��  G   ��  G   ��  FX  ��  FX      H   ,  �t  FX  �t  G   �<  G   �<  FX  �t  FX      H   ,  �  E�  �  FX  ��  FX  ��  E�  �  E�      H   ,  ��  A�  ��  Bp  ��  Bp  ��  A�  ��  A�      H   ,  �T  E�  �T  FX  �  FX  �  E�  �T  E�      H   ,  ��  G   ��  G�  �T  G�  �T  G   ��  G       H   ,  �  Bp  �  C8  ��  C8  ��  Bp  �  Bp      H   ,  ��  D   ��  D�  ��  D�  ��  D   ��  D       H   ,  �<  C8  �<  D   �  D   �  C8  �<  C8      H   ,  �  D   �  D�  ��  D�  ��  D   �  D       H   ,  �\  G�  �\  H�  �$  H�  �$  G�  �\  G�      H   ,  �  M`  �  N(  ��  N(  ��  M`  �  M`      H   ,  �  C8  �  D   ��  D   ��  C8  �  C8      H   ,  �D  G�  �D  H�  �  H�  �  G�  �D  G�      H   ,  �  Bp  �  C8  ��  C8  ��  Bp  �  Bp      H   ,  �  L�  �  M`  ��  M`  ��  L�  �  L�      H   ,  �  FX  �  G   ��  G   ��  FX  �  FX      H   ,  ��  G�  ��  H�  ͼ  H�  ͼ  G�  ��  G�      H   ,  �  K�  �  L�  ��  L�  ��  K�  �  K�      H   ,  ʜ  G�  ʜ  H�  �d  H�  �d  G�  ʜ  G�      H   ,  ��  G�  ��  H�  ƴ  H�  ƴ  G�  ��  G�      H   ,  �|  G�  �|  H�  �D  H�  �D  G�  �|  G�      H   ,  ƴ  G�  ƴ  H�  �|  H�  �|  G�  ƴ  G�      H   ,  �  E�  �  FX  ��  FX  ��  E�  �  E�      H   ,  ��  G�  ��  H�  Ô  H�  Ô  G�  ��  G�      H   ,  �  K  �  K�  ��  K�  ��  K  �  K      H   ,  �,  G�  �,  H�  ��  H�  ��  G�  �,  G�      H   ,  ��  G�  ��  H�  ʜ  H�  ʜ  G�  ��  G�      H   ,  �  N(  �  N�  ��  N�  ��  N(  �  N(      H   ,  �  J@  �  K  ��  K  ��  J@  �  J@      H   ,  Ô  G�  Ô  H�  �\  H�  �\  G�  Ô  G�      H   ,  �d  G�  �d  H�  �,  H�  �,  G�  �d  G�      H   ,  �  Ix  �  J@  ��  J@  ��  Ix  �  Ix      H   ,  �$  G�  �$  H�  ��  H�  ��  G�  �$  G�      H   ,  �  G�  �  H�  ��  H�  ��  G�  �  G�      H   ,  �  D�  �  E�  ��  E�  ��  D�  �  D�      H   ,  �  G   �  G�  ��  G�  ��  G   �  G       H   ,  �  H�  �  Ix  ��  Ix  ��  H�  �  H�      H   ,  ��  K  ��  K�  ʜ  K�  ʜ  K  ��  K      H   ,  �d  Ix  �d  J@  �,  J@  �,  Ix  �d  Ix      H   ,  ��  L�  ��  M`  ʜ  M`  ʜ  L�  ��  L�      H   ,  ʜ  L�  ʜ  M`  �d  M`  �d  L�  ʜ  L�      H   ,  ��  Ix  ��  J@  ʜ  J@  ʜ  Ix  ��  Ix      H   ,  �,  H�  �,  Ix  ��  Ix  ��  H�  �,  H�      H   ,  �d  H�  �d  Ix  �,  Ix  �,  H�  �d  H�      H   ,  ʜ  J@  ʜ  K  �d  K  �d  J@  ʜ  J@      H   ,  ʜ  K  ʜ  K�  �d  K�  �d  K  ʜ  K      H   ,  ��  K�  ��  L�  ʜ  L�  ʜ  K�  ��  K�      H   ,  ��  J@  ��  K  ʜ  K  ʜ  J@  ��  J@      H   ,  ��  M`  ��  N(  ʜ  N(  ʜ  M`  ��  M`      H   ,  ��  H�  ��  Ix  ʜ  Ix  ʜ  H�  ��  H�      H   ,  ʜ  H�  ʜ  Ix  �d  Ix  �d  H�  ʜ  H�      H   ,  ʜ  K�  ʜ  L�  �d  L�  �d  K�  ʜ  K�      H   ,  ʜ  Ix  ʜ  J@  �d  J@  �d  Ix  ʜ  Ix      H   ,  �\  K�  �\  L�  �$  L�  �$  K�  �\  K�      H   ,  ƴ  J@  ƴ  K  �|  K  �|  J@  ƴ  J@      H   ,  �|  K�  �|  L�  �D  L�  �D  K�  �|  K�      H   ,  ��  K  ��  K�  Ô  K�  Ô  K  ��  K      H   ,  Ô  L�  Ô  M`  �\  M`  �\  L�  Ô  L�      H   ,  ��  K  ��  K�  ƴ  K�  ƴ  K  ��  K      H   ,  ƴ  Ix  ƴ  J@  �|  J@  �|  Ix  ƴ  Ix      H   ,  ��  Ix  ��  J@  Ô  J@  Ô  Ix  ��  Ix      H   ,  �D  K  �D  K�  �  K�  �  K  �D  K      H   ,  ƴ  H�  ƴ  Ix  �|  Ix  �|  H�  ƴ  H�      H   ,  �|  J@  �|  K  �D  K  �D  J@  �|  J@      H   ,  ��  L�  ��  M`  ƴ  M`  ƴ  L�  ��  L�      H   ,  ��  N(  ��  N�  ƴ  N�  ƴ  N(  ��  N(      H   ,  Ô  K�  Ô  L�  �\  L�  �\  K�  Ô  K�      H   ,  �D  K�  �D  L�  �  L�  �  K�  �D  K�      H   ,  �\  K  �\  K�  �$  K�  �$  K  �\  K      H   ,  �$  N(  �$  N�  ��  N�  ��  N(  �$  N(      H   ,  Ô  K  Ô  K�  �\  K�  �\  K  Ô  K      H   ,  ��  J@  ��  K  ƴ  K  ƴ  J@  ��  J@      H   ,  ��  M`  ��  N(  ƴ  N(  ƴ  M`  ��  M`      H   ,  �$  M`  �$  N(  ��  N(  ��  M`  �$  M`      H   ,  �D  H�  �D  Ix  �  Ix  �  H�  �D  H�      H   ,  ƴ  N(  ƴ  N�  �|  N�  �|  N(  ƴ  N(      H   ,  Ô  J@  Ô  K  �\  K  �\  J@  Ô  J@      H   ,  �D  N(  �D  N�  �  N�  �  N(  �D  N(      H   ,  �$  L�  �$  M`  ��  M`  ��  L�  �$  L�      H   ,  �D  M`  �D  N(  �  N(  �  M`  �D  M`      H   ,  Ô  Ix  Ô  J@  �\  J@  �\  Ix  Ô  Ix      H   ,  �$  K�  �$  L�  ��  L�  ��  K�  �$  K�      H   ,  �\  L�  �\  M`  �$  M`  �$  L�  �\  L�      H   ,  Ô  N(  Ô  N�  �\  N�  �\  N(  Ô  N(      H   ,  Ô  H�  Ô  Ix  �\  Ix  �\  H�  Ô  H�      H   ,  ƴ  M`  ƴ  N(  �|  N(  �|  M`  ƴ  M`      H   ,  �$  K  �$  K�  ��  K�  ��  K  �$  K      H   ,  �\  N(  �\  N�  �$  N�  �$  N(  �\  N(      H   ,  �D  J@  �D  K  �  K  �  J@  �D  J@      H   ,  ƴ  L�  ƴ  M`  �|  M`  �|  L�  ƴ  L�      H   ,  ��  Ix  ��  J@  ƴ  J@  ƴ  Ix  ��  Ix      H   ,  �$  J@  �$  K  ��  K  ��  J@  �$  J@      H   ,  ��  K�  ��  L�  ƴ  L�  ƴ  K�  ��  K�      H   ,  ��  N(  ��  N�  Ô  N�  Ô  N(  ��  N(      H   ,  �\  J@  �\  K  �$  K  �$  J@  �\  J@      H   ,  �$  Ix  �$  J@  ��  J@  ��  Ix  �$  Ix      H   ,  �\  M`  �\  N(  �$  N(  �$  M`  �\  M`      H   ,  �$  H�  �$  Ix  ��  Ix  ��  H�  �$  H�      H   ,  ƴ  K�  ƴ  L�  �|  L�  �|  K�  ƴ  K�      H   ,  ��  K�  ��  L�  Ô  L�  Ô  K�  ��  K�      H   ,  ��  M`  ��  N(  Ô  N(  Ô  M`  ��  M`      H   ,  Ô  M`  Ô  N(  �\  N(  �\  M`  Ô  M`      H   ,  �D  L�  �D  M`  �  M`  �  L�  �D  L�      H   ,  �D  Ix  �D  J@  �  J@  �  Ix  �D  Ix      H   ,  �|  H�  �|  Ix  �D  Ix  �D  H�  �|  H�      H   ,  ƴ  K  ƴ  K�  �|  K�  �|  K  ƴ  K      H   ,  ��  H�  ��  Ix  ƴ  Ix  ƴ  H�  ��  H�      H   ,  �\  Ix  �\  J@  �$  J@  �$  Ix  �\  Ix      H   ,  �\  H�  �\  Ix  �$  Ix  �$  H�  �\  H�      H   ,  ��  L�  ��  M`  Ô  M`  Ô  L�  ��  L�      H   ,  ��  H�  ��  Ix  Ô  Ix  Ô  H�  ��  H�      H   ,  �|  N(  �|  N�  �D  N�  �D  N(  �|  N(      H   ,  ��  J@  ��  K  Ô  K  Ô  J@  ��  J@      H   ,  �|  K  �|  K�  �D  K�  �D  K  �|  K      H   ,  �|  M`  �|  N(  �D  N(  �D  M`  �|  M`      H   ,  �|  Ix  �|  J@  �D  J@  �D  Ix  �|  Ix      H   ,  �|  L�  �|  M`  �D  M`  �D  L�  �|  L�      H   ,  ��  D�  ��  E�  ƴ  E�  ƴ  D�  ��  D�      H   ,  ƴ  D   ƴ  D�  �|  D�  �|  D   ƴ  D       H   ,  �D  C8  �D  D   �  D   �  C8  �D  C8      H   ,  �\  A�  �\  Bp  �$  Bp  �$  A�  �\  A�      H   ,  �$  D   �$  D�  ��  D�  ��  D   �$  D       H   ,  ��  D�  ��  E�  Ô  E�  Ô  D�  ��  D�      H   ,  ��  Bp  ��  C8  Ô  C8  Ô  Bp  ��  Bp      H   ,  ƴ  C8  ƴ  D   �|  D   �|  C8  ƴ  C8      H   ,  �D  D   �D  D�  �  D�  �  D   �D  D       H   ,  �|  D   �|  D�  �D  D�  �D  D   �|  D       H   ,  �|  A�  �|  Bp  �D  Bp  �D  A�  �|  A�      H   ,  �$  D�  �$  E�  ��  E�  ��  D�  �$  D�      H   ,  �$  Bp  �$  C8  ��  C8  ��  Bp  �$  Bp      H   ,  �\  D   �\  D�  �$  D�  �$  D   �\  D       H   ,  ƴ  Bp  ƴ  C8  �|  C8  �|  Bp  ƴ  Bp      H   ,  ��  D   ��  D�  ƴ  D�  ƴ  D   ��  D       H   ,  Ô  Bp  Ô  C8  �\  C8  �\  Bp  Ô  Bp      H   ,  Ô  C8  Ô  D   �\  D   �\  C8  Ô  C8      H   ,  ��  G   ��  G�  ƴ  G�  ƴ  G   ��  G       H   ,  �\  FX  �\  G   �$  G   �$  FX  �\  FX      H   ,  ƴ  A�  ƴ  Bp  �|  Bp  �|  A�  ƴ  A�      H   ,  ��  D   ��  D�  Ô  D�  Ô  D   ��  D       H   ,  �|  D�  �|  E�  �D  E�  �D  D�  �|  D�      H   ,  �|  Bp  �|  C8  �D  C8  �D  Bp  �|  Bp      H   ,  ��  C8  ��  D   Ô  D   Ô  C8  ��  C8      H   ,  �D  G   �D  G�  �  G�  �  G   �D  G       H   ,  ��  C8  ��  D   ƴ  D   ƴ  C8  ��  C8      H   ,  Ô  G   Ô  G�  �\  G�  �\  G   Ô  G       H   ,  ƴ  G   ƴ  G�  �|  G�  �|  G   ƴ  G       H   ,  �|  E�  �|  FX  �D  FX  �D  E�  �|  E�      H   ,  ��  FX  ��  G   ƴ  G   ƴ  FX  ��  FX      H   ,  �|  C8  �|  D   �D  D   �D  C8  �|  C8      H   ,  �|  FX  �|  G   �D  G   �D  FX  �|  FX      H   ,  ��  E�  ��  FX  Ô  FX  Ô  E�  ��  E�      H   ,  ��  G   ��  G�  Ô  G�  Ô  G   ��  G       H   ,  ��  Bp  ��  C8  ƴ  C8  ƴ  Bp  ��  Bp      H   ,  �\  C8  �\  D   �$  D   �$  C8  �\  C8      H   ,  Ô  FX  Ô  G   �\  G   �\  FX  Ô  FX      H   ,  Ô  D   Ô  D�  �\  D�  �\  D   Ô  D       H   ,  ƴ  FX  ƴ  G   �|  G   �|  FX  ƴ  FX      H   ,  ��  E�  ��  FX  ƴ  FX  ƴ  E�  ��  E�      H   ,  �$  G   �$  G�  ��  G�  ��  G   �$  G       H   ,  �$  C8  �$  D   ��  D   ��  C8  �$  C8      H   ,  �D  A�  �D  Bp  �  Bp  �  A�  �D  A�      H   ,  �\  G   �\  G�  �$  G�  �$  G   �\  G       H   ,  ��  A�  ��  Bp  ƴ  Bp  ƴ  A�  ��  A�      H   ,  Ô  E�  Ô  FX  �\  FX  �\  E�  Ô  E�      H   ,  �$  FX  �$  G   ��  G   ��  FX  �$  FX      H   ,  �$  A�  �$  Bp  ��  Bp  ��  A�  �$  A�      H   ,  ƴ  E�  ƴ  FX  �|  FX  �|  E�  ƴ  E�      H   ,  �\  E�  �\  FX  �$  FX  �$  E�  �\  E�      H   ,  ��  A�  ��  Bp  Ô  Bp  Ô  A�  ��  A�      H   ,  �D  D�  �D  E�  �  E�  �  D�  �D  D�      H   ,  �D  Bp  �D  C8  �  C8  �  Bp  �D  Bp      H   ,  �\  Bp  �\  C8  �$  C8  �$  Bp  �\  Bp      H   ,  �|  G   �|  G�  �D  G�  �D  G   �|  G       H   ,  ƴ  D�  ƴ  E�  �|  E�  �|  D�  ƴ  D�      H   ,  �$  E�  �$  FX  ��  FX  ��  E�  �$  E�      H   ,  Ô  A�  Ô  Bp  �\  Bp  �\  A�  Ô  A�      H   ,  �D  FX  �D  G   �  G   �  FX  �D  FX      H   ,  �D  E�  �D  FX  �  FX  �  E�  �D  E�      H   ,  ��  FX  ��  G   Ô  G   Ô  FX  ��  FX      H   ,  Ô  D�  Ô  E�  �\  E�  �\  D�  Ô  D�      H   ,  �\  D�  �\  E�  �$  E�  �$  D�  �\  D�      H   ,  ��  D�  ��  E�  ͼ  E�  ͼ  D�  ��  D�      H   ,  �L  D   �L  D�  �  D�  �  D   �L  D       H   ,  �,  A�  �,  Bp  ��  Bp  ��  A�  �,  A�      H   ,  ΄  A�  ΄  Bp  �L  Bp  �L  A�  ΄  A�      H   ,  ��  D   ��  D�  ʜ  D�  ʜ  D   ��  D       H   ,  ͼ  FX  ͼ  G   ΄  G   ΄  FX  ͼ  FX      H   ,  ʜ  E�  ʜ  FX  �d  FX  �d  E�  ʜ  E�      H   ,  ʜ  G   ʜ  G�  �d  G�  �d  G   ʜ  G       H   ,  �L  A�  �L  Bp  �  Bp  �  A�  �L  A�      H   ,  �,  D   �,  D�  ��  D�  ��  D   �,  D       H   ,  �,  E�  �,  FX  ��  FX  ��  E�  �,  E�      H   ,  ͼ  A�  ͼ  Bp  ΄  Bp  ΄  A�  ͼ  A�      H   ,  �,  C8  �,  D   ��  D   ��  C8  �,  C8      H   ,  ͼ  E�  ͼ  FX  ΄  FX  ΄  E�  ͼ  E�      H   ,  ��  D   ��  D�  ͼ  D�  ͼ  D   ��  D       H   ,  �d  G   �d  G�  �,  G�  �,  G   �d  G       H   ,  �d  D�  �d  E�  �,  E�  �,  D�  �d  D�      H   ,  ��  FX  ��  G   ʜ  G   ʜ  FX  ��  FX      H   ,  �,  D�  �,  E�  ��  E�  ��  D�  �,  D�      H   ,  �L  C8  �L  D   �  D   �  C8  �L  C8      H   ,  ��  FX  ��  G   ͼ  G   ͼ  FX  ��  FX      H   ,  ͼ  D�  ͼ  E�  ΄  E�  ΄  D�  ͼ  D�      H   ,  ʜ  D   ʜ  D�  �d  D�  �d  D   ʜ  D       H   ,  �,  G   �,  G�  ��  G�  ��  G   �,  G       H   ,  ͼ  Bp  ͼ  C8  ΄  C8  ΄  Bp  ͼ  Bp      H   ,  �,  Bp  �,  C8  ��  C8  ��  Bp  �,  Bp      H   ,  �d  D   �d  D�  �,  D�  �,  D   �d  D       H   ,  ΄  D�  ΄  E�  �L  E�  �L  D�  ΄  D�      H   ,  ΄  C8  ΄  D   �L  D   �L  C8  ΄  C8      H   ,  ��  C8  ��  D   ͼ  D   ͼ  C8  ��  C8      H   ,  �L  D�  �L  E�  �  E�  �  D�  �L  D�      H   ,  �,  FX  �,  G   ��  G   ��  FX  �,  FX      H   ,  ͼ  D   ͼ  D�  ΄  D�  ΄  D   ͼ  D       H   ,  �d  FX  �d  G   �,  G   �,  FX  �d  FX      H   ,  �L  Bp  �L  C8  �  C8  �  Bp  �L  Bp      H   ,  ΄  FX  ΄  G   �L  G   �L  FX  ΄  FX      H   ,  ��  Bp  ��  C8  ͼ  C8  ͼ  Bp  ��  Bp      H   ,  ΄  D   ΄  D�  �L  D�  �L  D   ΄  D       H   ,  ��  E�  ��  FX  ʜ  FX  ʜ  E�  ��  E�      H   ,  ΄  E�  ΄  FX  �L  FX  �L  E�  ΄  E�      H   ,  ʜ  D�  ʜ  E�  �d  E�  �d  D�  ʜ  D�      H   ,  ��  E�  ��  FX  ͼ  FX  ͼ  E�  ��  E�      H   ,  �d  E�  �d  FX  �,  FX  �,  E�  �d  E�      H   ,  ��  D�  ��  E�  ʜ  E�  ʜ  D�  ��  D�      H   ,  ͼ  C8  ͼ  D   ΄  D   ΄  C8  ͼ  C8      H   ,  ��  A�  ��  Bp  ͼ  Bp  ͼ  A�  ��  A�      H   ,  ��  G   ��  G�  ʜ  G�  ʜ  G   ��  G       H   ,  �d  C8  �d  D   �,  D   �,  C8  �d  C8      H   ,  ΄  Bp  ΄  C8  �L  C8  �L  Bp  ΄  Bp      H   ,  ʜ  FX  ʜ  G   �d  G   �d  FX  ʜ  FX      H   ,  ͼ  G   ͼ  G�  ΄  G�  ΄  G   ͼ  G       H   ,  ��  C8  ��  D   ʜ  D   ʜ  C8  ��  C8      H   ,  ��  G   ��  G�  ͼ  G�  ͼ  G   ��  G       H   ,  �  jH  �  k  ��  k  ��  jH  �  jH      H   ,  �<  jH  �<  k  �  k  �  jH  �<  jH      H   ,  ��  jH  ��  k  �\  k  �\  jH  ��  jH      H   ,  ��  jH  ��  k  �t  k  �t  jH  ��  jH      H   ,  �T  p�  �T  qP  �  qP  �  p�  �T  p�      H   ,  �T  o�  �T  p�  �  p�  �  o�  �T  o�      H   ,  �T  n�  �T  o�  �  o�  �  n�  �T  n�      H   ,  �T  n0  �T  n�  �  n�  �  n0  �T  n0      H   ,  �T  mh  �T  n0  �  n0  �  mh  �T  mh      H   ,  �T  l�  �T  mh  �  mh  �  l�  �T  l�      H   ,  �T  k�  �T  l�  �  l�  �  k�  �T  k�      H   ,  �T  k  �T  k�  �  k�  �  k  �T  k      H   ,  �T  jH  �T  k  �  k  �  jH  �T  jH      H   ,  �t  jH  �t  k  �<  k  �<  jH  �t  jH      H   ,  ��  jH  ��  k  ��  k  ��  jH  ��  jH      H   ,  �  jH  �  k  ��  k  ��  jH  �  jH      H   ,  ��  jH  ��  k  ��  k  ��  jH  ��  jH      H   ,  ��  k  ��  k�  �t  k�  �t  k  ��  k      H   ,  �  n0  �  n�  ��  n�  ��  n0  �  n0      H   ,  �  mh  �  n0  ��  n0  ��  mh  �  mh      H   ,  �  l�  �  mh  ��  mh  ��  l�  �  l�      H   ,  �  k�  �  l�  ��  l�  ��  k�  �  k�      H   ,  �  k  �  k�  ��  k�  ��  k  �  k      H   ,  �<  l�  �<  mh  �  mh  �  l�  �<  l�      H   ,  �  o�  �  p�  ��  p�  ��  o�  �  o�      H   ,  �<  k�  �<  l�  �  l�  �  k�  �<  k�      H   ,  ��  mh  ��  n0  �t  n0  �t  mh  ��  mh      H   ,  �<  k  �<  k�  �  k�  �  k  �<  k      H   ,  �t  mh  �t  n0  �<  n0  �<  mh  �t  mh      H   ,  ��  k  ��  k�  ��  k�  ��  k  ��  k      H   ,  �t  l�  �t  mh  �<  mh  �<  l�  �t  l�      H   ,  �t  k�  �t  l�  �<  l�  �<  k�  �t  k�      H   ,  �t  k  �t  k�  �<  k�  �<  k  �t  k      H   ,  ��  n0  ��  n�  �t  n�  �t  n0  ��  n0      H   ,  ��  l�  ��  mh  �t  mh  �t  l�  ��  l�      H   ,  �  k�  �  l�  ��  l�  ��  k�  �  k�      H   ,  �  k  �  k�  ��  k�  ��  k  �  k      H   ,  ��  n�  ��  o�  ��  o�  ��  n�  ��  n�      H   ,  �  n�  �  o�  ��  o�  ��  n�  �  n�      H   ,  ��  n0  ��  n�  ��  n�  ��  n0  ��  n0      H   ,  ��  mh  ��  n0  ��  n0  ��  mh  ��  mh      H   ,  ��  l�  ��  mh  ��  mh  ��  l�  ��  l�      H   ,  ��  k�  ��  l�  ��  l�  ��  k�  ��  k�      H   ,  ��  k  ��  k�  ��  k�  ��  k  ��  k      H   ,  ��  k�  ��  l�  �t  l�  �t  k�  ��  k�      H   ,  ��  qP  ��  r  �T  r  �T  qP  ��  qP      H   ,  ��  qP  ��  r  ��  r  ��  qP  ��  qP      H   ,  �  qP  �  r  ��  r  ��  qP  �  qP      H   ,  ��  qP  ��  r  ��  r  ��  qP  ��  qP      H   ,  �L  u8  �L  v   �  v   �  u8  �L  u8      H   ,  �L  tp  �L  u8  �  u8  �  tp  �L  tp      H   ,  ��  qP  ��  r  ��  r  ��  qP  ��  qP      H   ,  �L  s�  �L  tp  �  tp  �  s�  �L  s�      H   ,  �L  r�  �L  s�  �  s�  �  r�  �L  r�      H   ,  �L  r  �L  r�  �  r�  �  r  �L  r      H   ,  �L  qP  �L  r  �  r  �  qP  �L  qP      H   ,  �L  p�  �L  qP  �  qP  �  p�  �L  p�      H   ,  �4  qP  �4  r  ��  r  ��  qP  �4  qP      H   ,  ��  qP  ��  r  ��  r  ��  qP  ��  qP      H   ,  ��  qP  ��  r  ��  r  ��  qP  ��  qP      H   ,  ��  qP  ��  r  �l  r  �l  qP  ��  qP      H   ,  ��  qP  ��  r  �L  r  �L  qP  ��  qP      H   ,  �l  qP  �l  r  �4  r  �4  qP  �l  qP      H   ,  ��  tp  ��  u8  ��  u8  ��  tp  ��  tp      H   ,  ��  r  ��  r�  �l  r�  �l  r  ��  r      H   ,  �4  r  �4  r�  ��  r�  ��  r  �4  r      H   ,  ��  s�  ��  tp  ��  tp  ��  s�  ��  s�      H   ,  ��  r�  ��  s�  ��  s�  ��  r�  ��  r�      H   ,  �  s�  �  tp  ��  tp  ��  s�  �  s�      H   ,  �  r�  �  s�  ��  s�  ��  r�  �  r�      H   ,  ��  r  ��  r�  ��  r�  ��  r  ��  r      H   ,  �  r  �  r�  ��  r�  ��  r  �  r      H   ,  �  tp  �  u8  ��  u8  ��  tp  �  tp      H   ,  ��  r  ��  r�  ��  r�  ��  r  ��  r      H   ,  ��  r�  ��  s�  �l  s�  �l  r�  ��  r�      H   ,  �l  s�  �l  tp  �4  tp  �4  s�  �l  s�      H   ,  ��  s�  ��  tp  �l  tp  �l  s�  ��  s�      H   ,  �l  r�  �l  s�  �4  s�  �4  r�  �l  r�      H   ,  �l  r  �l  r�  �4  r�  �4  r  �l  r      H   ,  �4  r�  �4  s�  ��  s�  ��  r�  �4  r�      H   ,  �  u8  �  v   �d  v   �d  u8  �  u8      H   ,  ��  u8  ��  v   ��  v   ��  u8  ��  u8      H   ,  ��  tp  ��  u8  ��  u8  ��  tp  ��  tp      H   ,  �  tp  �  u8  �d  u8  �d  tp  �  tp      H   ,  ��  u8  ��  v   ��  v   ��  u8  ��  u8      H   ,  ��  tp  ��  u8  ��  u8  ��  tp  ��  tp      H   ,  ��  s�  ��  tp  ��  tp  ��  s�  ��  s�      H   ,  �  s�  �  tp  �d  tp  �d  s�  �  s�      H   ,  �d  u8  �d  v   �,  v   �,  u8  �d  u8      H   ,  ��  tp  ��  u8  �L  u8  �L  tp  ��  tp      H   ,  �  r�  �  s�  �d  s�  �d  r�  �  r�      H   ,  ��  r�  ��  s�  ��  s�  ��  r�  ��  r�      H   ,  �d  r�  �d  s�  �,  s�  �,  r�  �d  r�      H   ,  ��  r  ��  r�  ��  r�  ��  r  ��  r      H   ,  �  r  �  r�  �d  r�  �d  r  �  r      H   ,  �d  tp  �d  u8  �,  u8  �,  tp  �d  tp      H   ,  ��  r�  ��  s�  ��  s�  ��  r�  ��  r�      H   ,  ~  r  ~  r�  ~�  r�  ~�  r  ~  r      H   ,  ��  s�  ��  tp  �L  tp  �L  s�  ��  s�      H   ,  �d  r  �d  r�  �,  r�  �,  r  �d  r      H   ,  ��  r�  ��  s�  �L  s�  �L  r�  ��  r�      H   ,  ~�  v�  ~�  w�  �  w�  �  v�  ~�  v�      H   ,  ��  r  ��  r�  �L  r�  �L  r  ��  r      H   ,  ~�  v   ~�  v�  �  v�  �  v   ~�  v       H   ,  ��  s�  ��  tp  ��  tp  ��  s�  ��  s�      H   ,  ~�  u8  ~�  v   �  v   �  u8  ~�  u8      H   ,  ~  u8  ~  v   ~�  v   ~�  u8  ~  u8      H   ,  ~�  tp  ~�  u8  �  u8  �  tp  ~�  tp      H   ,  ~  tp  ~  u8  ~�  u8  ~�  tp  ~  tp      H   ,  �d  s�  �d  tp  �,  tp  �,  s�  �d  s�      H   ,  ~  s�  ~  tp  ~�  tp  ~�  s�  ~  s�      H   ,  ~�  s�  ~�  tp  �  tp  �  s�  ~�  s�      H   ,  ��  r  ��  r�  ��  r�  ��  r  ��  r      H   ,  �  v�  �  w�  �d  w�  �d  v�  �  v�      H   ,  �  v   �  v�  �d  v�  �d  v   �  v       H   ,  ~�  r�  ~�  s�  �  s�  �  r�  ~�  r�      H   ,  �d  v   �d  v�  �,  v�  �,  v   �d  v       H   ,  ~  r�  ~  s�  ~�  s�  ~�  r�  ~  r�      H   ,  ~�  r  ~�  r�  �  r�  �  r  ~�  r      H   ,  ��  u8  ��  v   �L  v   �L  u8  ��  u8      H   ,  �,  v   �,  v�  ��  v�  ��  v   �,  v       H   ,  �d  v�  �d  w�  �,  w�  �,  v�  �d  v�      H   ,  ~  v�  ~  w�  ~�  w�  ~�  v�  ~  v�      H   ,  �,  u8  �,  v   ��  v   ��  u8  �,  u8      H   ,  ��  v   ��  v�  ��  v�  ��  v   ��  v       H   ,  �,  tp  �,  u8  ��  u8  ��  tp  �,  tp      H   ,  �,  s�  �,  tp  ��  tp  ��  s�  �,  s�      H   ,  �,  r�  �,  s�  ��  s�  ��  r�  �,  r�      H   ,  �,  r  �,  r�  ��  r�  ��  r  �,  r      H   ,  ��  v   ��  v�  ��  v�  ��  v   ��  v       H   ,  ~  v   ~  v�  ~�  v�  ~�  v   ~  v       H   ,  ��  p�  ��  qP  �L  qP  �L  p�  ��  p�      H   ,  �  o�  �  p�  ��  p�  ��  o�  �  o�      H   ,  ��  l�  ��  mh  ��  mh  ��  l�  ��  l�      H   ,  ��  n0  ��  n�  ��  n�  ��  n0  ��  n0      H   ,  ��  k�  ��  l�  ��  l�  ��  k�  ��  k�      H   ,  ��  p�  ��  qP  ��  qP  ��  p�  ��  p�      H   ,  �l  o�  �l  p�  �4  p�  �4  o�  �l  o�      H   ,  �  p�  �  qP  ��  qP  ��  p�  �  p�      H   ,  ��  p�  ��  qP  �l  qP  �l  p�  ��  p�      H   ,  ��  l�  ��  mh  ��  mh  ��  l�  ��  l�      H   ,  ��  o�  ��  p�  ��  p�  ��  o�  ��  o�      H   ,  �l  n0  �l  n�  �4  n�  �4  n0  �l  n0      H   ,  ��  o�  ��  p�  �l  p�  �l  o�  ��  o�      H   ,  ��  p�  ��  qP  �T  qP  �T  p�  ��  p�      H   ,  ��  n�  ��  o�  �T  o�  �T  n�  ��  n�      H   ,  �l  n�  �l  o�  �4  o�  �4  n�  �l  n�      H   ,  ��  n0  ��  n�  �T  n�  �T  n0  ��  n0      H   ,  �4  p�  �4  qP  ��  qP  ��  p�  �4  p�      H   ,  ��  p�  ��  qP  ��  qP  ��  p�  ��  p�      H   ,  ��  mh  ��  n0  �T  n0  �T  mh  ��  mh      H   ,  ��  mh  ��  n0  ��  n0  ��  mh  ��  mh      H   ,  ��  o�  ��  p�  ��  p�  ��  o�  ��  o�      H   ,  ��  k�  ��  l�  �T  l�  �T  k�  ��  k�      H   ,  �4  o�  �4  p�  ��  p�  ��  o�  �4  o�      H   ,  ��  n�  ��  o�  ��  o�  ��  n�  ��  n�      H   ,  ��  n�  ��  o�  �l  o�  �l  n�  ��  n�      H   ,  ��  n0  ��  n�  �l  n�  �l  n0  ��  n0      H   ,  �4  n�  �4  o�  ��  o�  ��  n�  �4  n�      H   ,  ��  o�  ��  p�  �T  p�  �T  o�  ��  o�      H   ,  �4  n0  �4  n�  ��  n�  ��  n0  �4  n0      H   ,  ��  k  ��  k�  �T  k�  �T  k  ��  k      H   ,  ��  p�  ��  qP  ��  qP  ��  p�  ��  p�      H   ,  ��  o�  ��  p�  ��  p�  ��  o�  ��  o�      H   ,  ��  n�  ��  o�  ��  o�  ��  n�  ��  n�      H   ,  ��  n�  ��  o�  ��  o�  ��  n�  ��  n�      H   ,  �4  mh  �4  n0  ��  n0  ��  mh  �4  mh      H   ,  �l  p�  �l  qP  �4  qP  �4  p�  �l  p�      H   ,  ��  n0  ��  n�  ��  n�  ��  n0  ��  n0      H   ,  ��  l�  ��  mh  �T  mh  �T  l�  ��  l�      H   ,  ��  mh  ��  n0  ��  n0  ��  mh  ��  mh      H   ,  �  e�  �  f`  �d  f`  �d  e�  �  e�      H   ,  ~  _X  ~  `   ~�  `   ~�  _X  ~  _X      H   ,  �d  `�  �d  a�  �,  a�  �,  `�  �d  `�      H   ,  �d  c@  �d  d  �,  d  �,  c@  �d  c@      H   ,  �  d�  �  e�  �d  e�  �d  d�  �  d�      H   ,  ��  d  ��  d�  ��  d�  ��  d  ��  d      H   ,  ~�  bx  ~�  c@  �  c@  �  bx  ~�  bx      H   ,  �  d  �  d�  �d  d�  �d  d  �  d      H   ,  �  c@  �  d  �d  d  �d  c@  �  c@      H   ,  ��  c@  ��  d  ��  d  ��  c@  ��  c@      H   ,  �  bx  �  c@  �d  c@  �d  bx  �  bx      H   ,  �  a�  �  bx  �d  bx  �d  a�  �  a�      H   ,  ~  d  ~  d�  ~�  d�  ~�  d  ~  d      H   ,  ��  bx  ��  c@  ��  c@  ��  bx  ��  bx      H   ,  �  `�  �  a�  �d  a�  �d  `�  �  `�      H   ,  ~�  `�  ~�  a�  �  a�  �  `�  ~�  `�      H   ,  �d  `   �d  `�  �,  `�  �,  `   �d  `       H   ,  �  `   �  `�  �d  `�  �d  `   �  `       H   ,  ~�  ]�  ~�  ^�  �  ^�  �  ]�  ~�  ]�      H   ,  �,  `�  �,  a�  ��  a�  ��  `�  �,  `�      H   ,  �  _X  �  `   �d  `   �d  _X  �  _X      H   ,  ~  g�  ~  h�  ~�  h�  ~�  g�  ~  g�      H   ,  ~  c@  ~  d  ~�  d  ~�  c@  ~  c@      H   ,  �  ^�  �  _X  �d  _X  �d  ^�  �  ^�      H   ,  ��  a�  ��  bx  ��  bx  ��  a�  ��  a�      H   ,  ~  ^�  ~  _X  ~�  _X  ~�  ^�  ~  ^�      H   ,  �  ]�  �  ^�  �d  ^�  �d  ]�  �  ]�      H   ,  �d  bx  �d  c@  �,  c@  �,  bx  �d  bx      H   ,  ~�  ]   ~�  ]�  �  ]�  �  ]   ~�  ]       H   ,  �  ]   �  ]�  �d  ]�  �d  ]   �  ]       H   ,  ��  `�  ��  a�  ��  a�  ��  `�  ��  `�      H   ,  �d  _X  �d  `   �,  `   �,  _X  �d  _X      H   ,  ~  g(  ~  g�  ~�  g�  ~�  g(  ~  g(      H   ,  �,  `   �,  `�  ��  `�  ��  `   �,  `       H   ,  �,  _X  �,  `   ��  `   ��  _X  �,  _X      H   ,  ~  bx  ~  c@  ~�  c@  ~�  bx  ~  bx      H   ,  ��  `   ��  `�  ��  `�  ��  `   ��  `       H   ,  �d  f`  �d  g(  �,  g(  �,  f`  �d  f`      H   ,  �,  ^�  �,  _X  ��  _X  ��  ^�  �,  ^�      H   ,  �d  ^�  �d  _X  �,  _X  �,  ^�  �d  ^�      H   ,  �,  ]�  �,  ^�  ��  ^�  ��  ]�  �,  ]�      H   ,  ��  _X  ��  `   ��  `   ��  _X  ��  _X      H   ,  ~  a�  ~  bx  ~�  bx  ~�  a�  ~  a�      H   ,  �d  e�  �d  f`  �,  f`  �,  e�  �d  e�      H   ,  �,  d  �,  d�  ��  d�  ��  d  �,  d      H   ,  �,  ]   �,  ]�  ��  ]�  ��  ]   �,  ]       H   ,  ��  ^�  ��  _X  ��  _X  ��  ^�  ��  ^�      H   ,  �d  ]�  �d  ^�  �,  ^�  �,  ]�  �d  ]�      H   ,  ~  `�  ~  a�  ~�  a�  ~�  `�  ~  `�      H   ,  �d  d�  �d  e�  �,  e�  �,  d�  �d  d�      H   ,  ~  ]�  ~  ^�  ~�  ^�  ~�  ]�  ~  ]�      H   ,  �d  a�  �d  bx  �,  bx  �,  a�  �d  a�      H   ,  ~  f`  ~  g(  ~�  g(  ~�  f`  ~  f`      H   ,  �,  e�  �,  f`  ��  f`  ��  e�  �,  e�      H   ,  ��  ]�  ��  ^�  ��  ^�  ��  ]�  ��  ]�      H   ,  ~�  `   ~�  `�  �  `�  �  `   ~�  `       H   ,  �,  c@  �,  d  ��  d  ��  c@  �,  c@      H   ,  �d  ]   �d  ]�  �,  ]�  �,  ]   �d  ]       H   ,  ~  `   ~  `�  ~�  `�  ~�  `   ~  `       H   ,  ~�  g�  ~�  h�  �  h�  �  g�  ~�  g�      H   ,  ~�  g(  ~�  g�  �  g�  �  g(  ~�  g(      H   ,  �d  d  �d  d�  �,  d�  �,  d  �d  d      H   ,  ~�  a�  ~�  bx  �  bx  �  a�  ~�  a�      H   ,  ��  ]   ��  ]�  ��  ]�  ��  ]   ��  ]       H   ,  ~  e�  ~  f`  ~�  f`  ~�  e�  ~  e�      H   ,  ~�  f`  ~�  g(  �  g(  �  f`  ~�  f`      H   ,  �,  d�  �,  e�  ��  e�  ��  d�  �,  d�      H   ,  �  g(  �  g�  �d  g�  �d  g(  �  g(      H   ,  ~�  e�  ~�  f`  �  f`  �  e�  ~�  e�      H   ,  ~�  _X  ~�  `   �  `   �  _X  ~�  _X      H   ,  ~�  d�  ~�  e�  �  e�  �  d�  ~�  d�      H   ,  �,  bx  �,  c@  ��  c@  ��  bx  �,  bx      H   ,  ~�  d  ~�  d�  �  d�  �  d  ~�  d      H   ,  �  f`  �  g(  �d  g(  �d  f`  �  f`      H   ,  ~  d�  ~  e�  ~�  e�  ~�  d�  ~  d�      H   ,  ~�  c@  ~�  d  �  d  �  c@  ~�  c@      H   ,  ~�  ^�  ~�  _X  �  _X  �  ^�  ~�  ^�      H   ,  �,  a�  �,  bx  ��  bx  ��  a�  �,  a�      H   ,  ~  ]   ~  ]�  ~�  ]�  ~�  ]   ~  ]       H   ,  �\  c@  �\  d  �$  d  �$  c@  �\  c@      H   ,  �\  bx  �\  c@  �$  c@  �$  bx  �\  bx      H   ,  ��  c@  ��  d  ��  d  ��  c@  ��  c@      H   ,  �\  i�  �\  jH  �$  jH  �$  i�  �\  i�      H   ,  �\  h�  �\  i�  �$  i�  �$  h�  �\  h�      H   ,  �\  g�  �\  h�  �$  h�  �$  g�  �\  g�      H   ,  �\  g(  �\  g�  �$  g�  �$  g(  �\  g(      H   ,  �$  c@  �$  d  ��  d  ��  c@  �$  c@      H   ,  �D  c@  �D  d  �  d  �  c@  �D  c@      H   ,  ��  c@  ��  d  �\  d  �\  c@  ��  c@      H   ,  �\  f`  �\  g(  �$  g(  �$  f`  �\  f`      H   ,  �|  c@  �|  d  �D  d  �D  c@  �|  c@      H   ,  �\  e�  �\  f`  �$  f`  �$  e�  �\  e�      H   ,  �  c@  �  d  ��  d  ��  c@  �  c@      H   ,  �\  d�  �\  e�  �$  e�  �$  d�  �\  d�      H   ,  ��  c@  ��  d  �|  d  �|  c@  ��  c@      H   ,  �\  d  �\  d�  �$  d�  �$  d  �\  d      H   ,  �$  g(  �$  g�  ��  g�  ��  g(  �$  g(      H   ,  ��  g(  ��  g�  ��  g�  ��  g(  ��  g(      H   ,  �$  h�  �$  i�  ��  i�  ��  h�  �$  h�      H   ,  �|  e�  �|  f`  �D  f`  �D  e�  �|  e�      H   ,  ��  f`  ��  g(  �|  g(  �|  f`  ��  f`      H   ,  �|  d�  �|  e�  �D  e�  �D  d�  �|  d�      H   ,  ��  d  ��  d�  ��  d�  ��  d  ��  d      H   ,  ��  d�  ��  e�  ��  e�  ��  d�  ��  d�      H   ,  �$  f`  �$  g(  ��  g(  ��  f`  �$  f`      H   ,  �|  d  �|  d�  �D  d�  �D  d  �|  d      H   ,  �$  e�  �$  f`  ��  f`  ��  e�  �$  e�      H   ,  ��  e�  ��  f`  �|  f`  �|  e�  ��  e�      H   ,  ��  f`  ��  g(  ��  g(  ��  f`  ��  f`      H   ,  �$  g�  �$  h�  ��  h�  ��  g�  �$  g�      H   ,  ��  d�  ��  e�  �|  e�  �|  d�  ��  d�      H   ,  ��  e�  ��  f`  ��  f`  ��  e�  ��  e�      H   ,  �  d  �  d�  ��  d�  ��  d  �  d      H   ,  �$  d�  �$  e�  ��  e�  ��  d�  �$  d�      H   ,  ��  d  ��  d�  �|  d�  �|  d  ��  d      H   ,  �D  d�  �D  e�  �  e�  �  d�  �D  d�      H   ,  ��  g�  ��  h�  ��  h�  ��  g�  ��  g�      H   ,  �$  d  �$  d�  ��  d�  ��  d  �$  d      H   ,  �D  d  �D  d�  �  d�  �  d  �D  d      H   ,  ��  d  ��  d�  �\  d�  �\  d  ��  d      H   ,  �  g�  �  h�  ��  h�  ��  g�  �  g�      H   ,  �<  f`  �<  g(  �  g(  �  f`  �<  f`      H   ,  �  g(  �  g�  ��  g�  ��  g(  �  g(      H   ,  ��  g�  ��  h�  �\  h�  �\  g�  ��  g�      H   ,  ��  e�  ��  f`  �\  f`  �\  e�  ��  e�      H   ,  ��  h�  ��  i�  ��  i�  ��  h�  ��  h�      H   ,  �t  g(  �t  g�  �<  g�  �<  g(  �t  g(      H   ,  ��  i�  ��  jH  �\  jH  �\  i�  ��  i�      H   ,  �  f`  �  g(  ��  g(  ��  f`  �  f`      H   ,  �  e�  �  f`  ��  f`  ��  e�  �  e�      H   ,  ��  i�  ��  jH  ��  jH  ��  i�  ��  i�      H   ,  ��  i�  ��  jH  ��  jH  ��  i�  ��  i�      H   ,  ��  g(  ��  g�  ��  g�  ��  g(  ��  g(      H   ,  ��  d�  ��  e�  ��  e�  ��  d�  ��  d�      H   ,  ��  d�  ��  e�  �\  e�  �\  d�  ��  d�      H   ,  ��  h�  ��  i�  ��  i�  ��  h�  ��  h�      H   ,  �<  i�  �<  jH  �  jH  �  i�  �<  i�      H   ,  ��  g(  ��  g�  �\  g�  �\  g(  ��  g(      H   ,  ��  h�  ��  i�  �t  i�  �t  h�  ��  h�      H   ,  �<  h�  �<  i�  �  i�  �  h�  �<  h�      H   ,  ��  h�  ��  i�  �\  i�  �\  h�  ��  h�      H   ,  ��  g�  ��  h�  ��  h�  ��  g�  ��  g�      H   ,  �  i�  �  jH  ��  jH  ��  i�  �  i�      H   ,  ��  i�  ��  jH  �t  jH  �t  i�  ��  i�      H   ,  ��  f`  ��  g(  ��  g(  ��  f`  ��  f`      H   ,  �<  g�  �<  h�  �  h�  �  g�  �<  g�      H   ,  �t  g�  �t  h�  �<  h�  �<  g�  �t  g�      H   ,  �  i�  �  jH  ��  jH  ��  i�  �  i�      H   ,  ��  g�  ��  h�  �t  h�  �t  g�  ��  g�      H   ,  ��  e�  ��  f`  ��  f`  ��  e�  ��  e�      H   ,  �<  g(  �<  g�  �  g�  �  g(  �<  g(      H   ,  ��  d  ��  d�  ��  d�  ��  d  ��  d      H   ,  �t  i�  �t  jH  �<  jH  �<  i�  �t  i�      H   ,  �t  h�  �t  i�  �<  i�  �<  h�  �t  h�      H   ,  �  h�  �  i�  ��  i�  ��  h�  �  h�      H   ,  ��  f`  ��  g(  �\  g(  �\  f`  ��  f`      H   ,  ��  a�  ��  bx  ��  bx  ��  a�  ��  a�      H   ,  ��  bx  ��  c@  ��  c@  ��  bx  ��  bx      H   ,  ��  `   ��  `�  �d  `�  �d  `   ��  `       H   ,  ��  ]�  ��  ^�  ��  ^�  ��  ]�  ��  ]�      H   ,  ��  a�  ��  bx  �d  bx  �d  a�  ��  a�      H   ,  ��  `   ��  `�  �|  `�  �|  `   ��  `       H   ,  ��  ^�  ��  _X  �d  _X  �d  ^�  ��  ^�      H   ,  ��  `   ��  `�  ��  `�  ��  `   ��  `       H   ,  �D  bx  �D  c@  �  c@  �  bx  �D  bx      H   ,  �|  bx  �|  c@  �D  c@  �D  bx  �|  bx      H   ,  �D  `�  �D  a�  �  a�  �  `�  �D  `�      H   ,  �D  ]   �D  ]�  �  ]�  �  ]   �D  ]       H   ,  ��  ]   ��  ]�  �d  ]�  �d  ]   ��  ]       H   ,  ��  _X  ��  `   ��  `   ��  _X  ��  _X      H   ,  ��  ]   ��  ]�  ��  ]�  ��  ]   ��  ]       H   ,  �D  `   �D  `�  �  `�  �  `   �D  `       H   ,  �$  bx  �$  c@  ��  c@  ��  bx  �$  bx      H   ,  �|  a�  �|  bx  �D  bx  �D  a�  �|  a�      H   ,  ��  _X  ��  `   �|  `   �|  _X  ��  _X      H   ,  ��  a�  ��  bx  �|  bx  �|  a�  ��  a�      H   ,  ��  _X  ��  `   �d  `   �d  _X  ��  _X      H   ,  �D  _X  �D  `   �  `   �  _X  �D  _X      H   ,  ��  bx  ��  c@  �|  c@  �|  bx  ��  bx      H   ,  �|  `�  �|  a�  �D  a�  �D  `�  �|  `�      H   ,  ��  `�  ��  a�  �d  a�  �d  `�  ��  `�      H   ,  �  bx  �  c@  ��  c@  ��  bx  �  bx      H   ,  �  a�  �  bx  ��  bx  ��  a�  �  a�      H   ,  ��  `�  ��  a�  ��  a�  ��  `�  ��  `�      H   ,  �  `�  �  a�  ��  a�  ��  `�  �  `�      H   ,  ��  ^�  ��  _X  ��  _X  ��  ^�  ��  ^�      H   ,  �  `   �  `�  ��  `�  ��  `   �  `       H   ,  �|  `   �|  `�  �D  `�  �D  `   �|  `       H   ,  �  _X  �  `   ��  `   ��  _X  �  _X      H   ,  �  ^�  �  _X  ��  _X  ��  ^�  �  ^�      H   ,  ��  a�  ��  bx  ��  bx  ��  a�  ��  a�      H   ,  �  ]�  �  ^�  ��  ^�  ��  ]�  �  ]�      H   ,  �D  ^�  �D  _X  �  _X  �  ^�  �D  ^�      H   ,  �|  _X  �|  `   �D  `   �D  _X  �|  _X      H   ,  �  ]   �  ]�  ��  ]�  ��  ]   �  ]       H   ,  �D  ]�  �D  ^�  �  ^�  �  ]�  �D  ]�      H   ,  ��  `�  ��  a�  �|  a�  �|  `�  ��  `�      H   ,  ��  ]�  ��  ^�  �d  ^�  �d  ]�  ��  ]�      H   ,  �D  a�  �D  bx  �  bx  �  a�  �D  a�      H   ,  ��  `�  ��  a�  ��  a�  ��  `�  ��  `�      H   ,  �|  ^�  �|  _X  �D  _X  �D  ^�  �|  ^�      H   ,  ��  bx  ��  c@  ��  c@  ��  bx  ��  bx      H   ,  �$  a�  �$  bx  ��  bx  ��  a�  �$  a�      H   ,  {�  jH  {�  k  ||  k  ||  jH  {�  jH      H   ,  z�  jH  z�  k  {�  k  {�  jH  z�  jH      H   ,  w�  jH  w�  k  x�  k  x�  jH  w�  jH      H   ,  x�  jH  x�  k  y\  k  y\  jH  x�  jH      H   ,  y\  jH  y\  k  z$  k  z$  jH  y\  jH      H   ,  z$  jH  z$  k  z�  k  z�  jH  z$  jH      H   ,  z�  k  z�  k�  {�  k�  {�  k  z�  k      H   ,  {�  k  {�  k�  ||  k�  ||  k  {�  k      H   ,  {�  u8  {�  v   ||  v   ||  u8  {�  u8      H   ,  {�  n0  {�  n�  ||  n�  ||  n0  {�  n0      H   ,  x�  n0  x�  n�  y\  n�  y\  n0  x�  n0      H   ,  ||  tp  ||  u8  }D  u8  }D  tp  ||  tp      H   ,  x�  qP  x�  r  y\  r  y\  qP  x�  qP      H   ,  y\  s�  y\  tp  z$  tp  z$  s�  y\  s�      H   ,  {�  tp  {�  u8  ||  u8  ||  tp  {�  tp      H   ,  }D  v   }D  v�  ~  v�  ~  v   }D  v       H   ,  w�  o�  w�  p�  x�  p�  x�  o�  w�  o�      H   ,  z�  r  z�  r�  {�  r�  {�  r  z�  r      H   ,  }D  u8  }D  v   ~  v   ~  u8  }D  u8      H   ,  y\  r�  y\  s�  z$  s�  z$  r�  y\  r�      H   ,  }D  tp  }D  u8  ~  u8  ~  tp  }D  tp      H   ,  x�  mh  x�  n0  y\  n0  y\  mh  x�  mh      H   ,  w�  n�  w�  o�  x�  o�  x�  n�  w�  n�      H   ,  }D  s�  }D  tp  ~  tp  ~  s�  }D  s�      H   ,  ||  s�  ||  tp  }D  tp  }D  s�  ||  s�      H   ,  y\  r  y\  r�  z$  r�  z$  r  y\  r      H   ,  {�  v   {�  v�  ||  v�  ||  v   {�  v       H   ,  }D  r�  }D  s�  ~  s�  ~  r�  }D  r�      H   ,  z�  n0  z�  n�  {�  n�  {�  n0  z�  n0      H   ,  z�  tp  z�  u8  {�  u8  {�  tp  z�  tp      H   ,  }D  r  }D  r�  ~  r�  ~  r  }D  r      H   ,  y\  qP  y\  r  z$  r  z$  qP  y\  qP      H   ,  }D  qP  }D  r  ~  r  ~  qP  }D  qP      H   ,  w�  n0  w�  n�  x�  n�  x�  n0  w�  n0      H   ,  {�  s�  {�  tp  ||  tp  ||  s�  {�  s�      H   ,  y\  p�  y\  qP  z$  qP  z$  p�  y\  p�      H   ,  x�  l�  x�  mh  y\  mh  y\  l�  x�  l�      H   ,  ||  r�  ||  s�  }D  s�  }D  r�  ||  r�      H   ,  w�  mh  w�  n0  x�  n0  x�  mh  w�  mh      H   ,  z�  l�  z�  mh  {�  mh  {�  l�  z�  l�      H   ,  y\  o�  y\  p�  z$  p�  z$  o�  y\  o�      H   ,  z�  qP  z�  r  {�  r  {�  qP  z�  qP      H   ,  y\  n�  y\  o�  z$  o�  z$  n�  y\  n�      H   ,  x�  k�  x�  l�  y\  l�  y\  k�  x�  k�      H   ,  w�  l�  w�  mh  x�  mh  x�  l�  w�  l�      H   ,  ||  r  ||  r�  }D  r�  }D  r  ||  r      H   ,  y\  n0  y\  n�  z$  n�  z$  n0  y\  n0      H   ,  x�  p�  x�  qP  y\  qP  y\  p�  x�  p�      H   ,  w�  k�  w�  l�  x�  l�  x�  k�  w�  k�      H   ,  {�  r�  {�  s�  ||  s�  ||  r�  {�  r�      H   ,  y\  mh  y\  n0  z$  n0  z$  mh  y\  mh      H   ,  x�  k  x�  k�  y\  k�  y\  k  x�  k      H   ,  w�  k  w�  k�  x�  k�  x�  k  w�  k      H   ,  y\  l�  y\  mh  z$  mh  z$  l�  y\  l�      H   ,  ||  qP  ||  r  }D  r  }D  qP  ||  qP      H   ,  z$  tp  z$  u8  z�  u8  z�  tp  z$  tp      H   ,  x�  r  x�  r�  y\  r�  y\  r  x�  r      H   ,  y\  k�  y\  l�  z$  l�  z$  k�  y\  k�      H   ,  z$  s�  z$  tp  z�  tp  z�  s�  z$  s�      H   ,  {�  r  {�  r�  ||  r�  ||  r  {�  r      H   ,  {�  mh  {�  n0  ||  n0  ||  mh  {�  mh      H   ,  z�  u8  z�  v   {�  v   {�  u8  z�  u8      H   ,  z$  r�  z$  s�  z�  s�  z�  r�  z$  r�      H   ,  z�  s�  z�  tp  {�  tp  {�  s�  z�  s�      H   ,  y\  k  y\  k�  z$  k�  z$  k  y\  k      H   ,  z�  p�  z�  qP  {�  qP  {�  p�  z�  p�      H   ,  ||  p�  ||  qP  }D  qP  }D  p�  ||  p�      H   ,  z$  r  z$  r�  z�  r�  z�  r  z$  r      H   ,  {�  l�  {�  mh  ||  mh  ||  l�  {�  l�      H   ,  x�  o�  x�  p�  y\  p�  y\  o�  x�  o�      H   ,  z$  qP  z$  r  z�  r  z�  qP  z$  qP      H   ,  z�  k�  z�  l�  {�  l�  {�  k�  z�  k�      H   ,  z$  p�  z$  qP  z�  qP  z�  p�  z$  p�      H   ,  z$  o�  z$  p�  z�  p�  z�  o�  z$  o�      H   ,  z$  n�  z$  o�  z�  o�  z�  n�  z$  n�      H   ,  z$  n0  z$  n�  z�  n�  z�  n0  z$  n0      H   ,  {�  qP  {�  r  ||  r  ||  qP  {�  qP      H   ,  ||  v   ||  v�  }D  v�  }D  v   ||  v       H   ,  z$  mh  z$  n0  z�  n0  z�  mh  z$  mh      H   ,  z$  l�  z$  mh  z�  mh  z�  l�  z$  l�      H   ,  z�  o�  z�  p�  {�  p�  {�  o�  z�  o�      H   ,  z$  k�  z$  l�  z�  l�  z�  k�  z$  k�      H   ,  {�  p�  {�  qP  ||  qP  ||  p�  {�  p�      H   ,  z�  mh  z�  n0  {�  n0  {�  mh  z�  mh      H   ,  z$  k  z$  k�  z�  k�  z�  k  z$  k      H   ,  {�  k�  {�  l�  ||  l�  ||  k�  {�  k�      H   ,  {�  o�  {�  p�  ||  p�  ||  o�  {�  o�      H   ,  x�  n�  x�  o�  y\  o�  y\  n�  x�  n�      H   ,  {�  n�  {�  o�  ||  o�  ||  n�  {�  n�      H   ,  z�  r�  z�  s�  {�  s�  {�  r�  z�  r�      H   ,  ||  u8  ||  v   }D  v   }D  u8  ||  u8      H   ,  z�  n�  z�  o�  {�  o�  {�  n�  z�  n�      H   ,  x�  c@  x�  d  y\  d  y\  c@  x�  c@      H   ,  w  d  w  d�  w�  d�  w�  d  w  d      H   ,  w  _X  w  `   w�  `   w�  _X  w  _X      H   ,  w�  c@  w�  d  x�  d  x�  c@  w�  c@      H   ,  s�  c@  s�  d  t�  d  t�  c@  s�  c@      H   ,  w  `   w  `�  w�  `�  w�  `   w  `       H   ,  w  ^�  w  _X  w�  _X  w�  ^�  w  ^�      H   ,  }D  c@  }D  d  ~  d  ~  c@  }D  c@      H   ,  w  a�  w  bx  w�  bx  w�  a�  w  a�      H   ,  w  c@  w  d  w�  d  w�  c@  w  c@      H   ,  w  ]�  w  ^�  w�  ^�  w�  ]�  w  ]�      H   ,  t�  c@  t�  d  ut  d  ut  c@  t�  c@      H   ,  z�  c@  z�  d  {�  d  {�  c@  z�  c@      H   ,  ut  c@  ut  d  v<  d  v<  c@  ut  c@      H   ,  y\  c@  y\  d  z$  d  z$  c@  y\  c@      H   ,  v<  c@  v<  d  w  d  w  c@  v<  c@      H   ,  w  ]   w  ]�  w�  ]�  w�  ]   w  ]       H   ,  {�  c@  {�  d  ||  d  ||  c@  {�  c@      H   ,  w  g�  w  h�  w�  h�  w�  g�  w  g�      H   ,  w  g(  w  g�  w�  g�  w�  g(  w  g(      H   ,  w  d�  w  e�  w�  e�  w�  d�  w  d�      H   ,  ||  c@  ||  d  }D  d  }D  c@  ||  c@      H   ,  w  f`  w  g(  w�  g(  w�  f`  w  f`      H   ,  w  `�  w  a�  w�  a�  w�  `�  w  `�      H   ,  w  bx  w  c@  w�  c@  w�  bx  w  bx      H   ,  w  e�  w  f`  w�  f`  w�  e�  w  e�      H   ,  z$  c@  z$  d  z�  d  z�  c@  z$  c@      H   ,  {�  f`  {�  g(  ||  g(  ||  f`  {�  f`      H   ,  x�  d�  x�  e�  y\  e�  y\  d�  x�  d�      H   ,  }D  h�  }D  i�  ~  i�  ~  h�  }D  h�      H   ,  {�  g(  {�  g�  ||  g�  ||  g(  {�  g(      H   ,  {�  d  {�  d�  ||  d�  ||  d  {�  d      H   ,  x�  e�  x�  f`  y\  f`  y\  e�  x�  e�      H   ,  }D  d�  }D  e�  ~  e�  ~  d�  }D  d�      H   ,  }D  g�  }D  h�  ~  h�  ~  g�  }D  g�      H   ,  ||  d  ||  d�  }D  d�  }D  d  ||  d      H   ,  w�  d  w�  d�  x�  d�  x�  d  w�  d      H   ,  }D  d  }D  d�  ~  d�  ~  d  }D  d      H   ,  {�  h�  {�  i�  ||  i�  ||  h�  {�  h�      H   ,  z�  i�  z�  jH  {�  jH  {�  i�  z�  i�      H   ,  w�  i�  w�  jH  x�  jH  x�  i�  w�  i�      H   ,  z�  f`  z�  g(  {�  g(  {�  f`  z�  f`      H   ,  z�  g(  z�  g�  {�  g�  {�  g(  z�  g(      H   ,  z�  e�  z�  f`  {�  f`  {�  e�  z�  e�      H   ,  w�  h�  w�  i�  x�  i�  x�  h�  w�  h�      H   ,  y\  i�  y\  jH  z$  jH  z$  i�  y\  i�      H   ,  x�  i�  x�  jH  y\  jH  y\  i�  x�  i�      H   ,  ||  h�  ||  i�  }D  i�  }D  h�  ||  h�      H   ,  x�  d  x�  d�  y\  d�  y\  d  x�  d      H   ,  w�  g�  w�  h�  x�  h�  x�  g�  w�  g�      H   ,  y\  h�  y\  i�  z$  i�  z$  h�  y\  h�      H   ,  {�  e�  {�  f`  ||  f`  ||  e�  {�  e�      H   ,  z�  d  z�  d�  {�  d�  {�  d  z�  d      H   ,  w�  g(  w�  g�  x�  g�  x�  g(  w�  g(      H   ,  y\  g�  y\  h�  z$  h�  z$  g�  y\  g�      H   ,  x�  h�  x�  i�  y\  i�  y\  h�  x�  h�      H   ,  ||  g�  ||  h�  }D  h�  }D  g�  ||  g�      H   ,  y\  g(  y\  g�  z$  g�  z$  g(  y\  g(      H   ,  }D  g(  }D  g�  ~  g�  ~  g(  }D  g(      H   ,  {�  g�  {�  h�  ||  h�  ||  g�  {�  g�      H   ,  {�  i�  {�  jH  ||  jH  ||  i�  {�  i�      H   ,  ||  d�  ||  e�  }D  e�  }D  d�  ||  d�      H   ,  w�  f`  w�  g(  x�  g(  x�  f`  w�  f`      H   ,  z�  h�  z�  i�  {�  i�  {�  h�  z�  h�      H   ,  z$  i�  z$  jH  z�  jH  z�  i�  z$  i�      H   ,  y\  f`  y\  g(  z$  g(  z$  f`  y\  f`      H   ,  z�  d�  z�  e�  {�  e�  {�  d�  z�  d�      H   ,  x�  g�  x�  h�  y\  h�  y\  g�  x�  g�      H   ,  z$  h�  z$  i�  z�  i�  z�  h�  z$  h�      H   ,  ||  g(  ||  g�  }D  g�  }D  g(  ||  g(      H   ,  z$  g�  z$  h�  z�  h�  z�  g�  z$  g�      H   ,  }D  f`  }D  g(  ~  g(  ~  f`  }D  f`      H   ,  y\  e�  y\  f`  z$  f`  z$  e�  y\  e�      H   ,  z$  g(  z$  g�  z�  g�  z�  g(  z$  g(      H   ,  z$  f`  z$  g(  z�  g(  z�  f`  z$  f`      H   ,  w�  e�  w�  f`  x�  f`  x�  e�  w�  e�      H   ,  z$  e�  z$  f`  z�  f`  z�  e�  z$  e�      H   ,  z$  d�  z$  e�  z�  e�  z�  d�  z$  d�      H   ,  y\  d�  y\  e�  z$  e�  z$  d�  y\  d�      H   ,  {�  d�  {�  e�  ||  e�  ||  d�  {�  d�      H   ,  x�  g(  x�  g�  y\  g�  y\  g(  x�  g(      H   ,  z$  d  z$  d�  z�  d�  z�  d  z$  d      H   ,  ||  f`  ||  g(  }D  g(  }D  f`  ||  f`      H   ,  }D  e�  }D  f`  ~  f`  ~  e�  }D  e�      H   ,  y\  d  y\  d�  z$  d�  z$  d  y\  d      H   ,  x�  f`  x�  g(  y\  g(  y\  f`  x�  f`      H   ,  z�  g�  z�  h�  {�  h�  {�  g�  z�  g�      H   ,  ||  e�  ||  f`  }D  f`  }D  e�  ||  e�      H   ,  w�  d�  w�  e�  x�  e�  x�  d�  w�  d�      H   ,  v<  d�  v<  e�  w  e�  w  d�  v<  d�      H   ,  t�  d  t�  d�  ut  d�  ut  d  t�  d      H   ,  v<  e�  v<  f`  w  f`  w  e�  v<  e�      H   ,  ut  f`  ut  g(  v<  g(  v<  f`  ut  f`      H   ,  t�  e�  t�  f`  ut  f`  ut  e�  t�  e�      H   ,  s�  d  s�  d�  t�  d�  t�  d  s�  d      H   ,  ut  e�  ut  f`  v<  f`  v<  e�  ut  e�      H   ,  v<  d  v<  d�  w  d�  w  d  v<  d      H   ,  ut  d�  ut  e�  v<  e�  v<  d�  ut  d�      H   ,  ut  d  ut  d�  v<  d�  v<  d  ut  d      H   ,  t�  d�  t�  e�  ut  e�  ut  d�  t�  d�      H   ,  v<  g(  v<  g�  w  g�  w  g(  v<  g(      H   ,  v<  f`  v<  g(  w  g(  w  f`  v<  f`      H   ,  t�  bx  t�  c@  ut  c@  ut  bx  t�  bx      H   ,  t�  ]   t�  ]�  ut  ]�  ut  ]   t�  ]       H   ,  ut  `�  ut  a�  v<  a�  v<  `�  ut  `�      H   ,  ut  ]�  ut  ^�  v<  ^�  v<  ]�  ut  ]�      H   ,  s�  `   s�  `�  t�  `�  t�  `   s�  `       H   ,  s�  bx  s�  c@  t�  c@  t�  bx  s�  bx      H   ,  s�  ]   s�  ]�  t�  ]�  t�  ]   s�  ]       H   ,  v<  bx  v<  c@  w  c@  w  bx  v<  bx      H   ,  v<  ]   v<  ]�  w  ]�  w  ]   v<  ]       H   ,  ut  `   ut  `�  v<  `�  v<  `   ut  `       H   ,  t�  `   t�  `�  ut  `�  ut  `   t�  `       H   ,  s�  a�  s�  bx  t�  bx  t�  a�  s�  a�      H   ,  ut  bx  ut  c@  v<  c@  v<  bx  ut  bx      H   ,  t�  a�  t�  bx  ut  bx  ut  a�  t�  a�      H   ,  ut  ^�  ut  _X  v<  _X  v<  ^�  ut  ^�      H   ,  s�  _X  s�  `   t�  `   t�  _X  s�  _X      H   ,  ut  a�  ut  bx  v<  bx  v<  a�  ut  a�      H   ,  t�  _X  t�  `   ut  `   ut  _X  t�  _X      H   ,  s�  ]�  s�  ^�  t�  ^�  t�  ]�  s�  ]�      H   ,  ut  ]   ut  ]�  v<  ]�  v<  ]   ut  ]       H   ,  v<  _X  v<  `   w  `   w  _X  v<  _X      H   ,  v<  ]�  v<  ^�  w  ^�  w  ]�  v<  ]�      H   ,  t�  ^�  t�  _X  ut  _X  ut  ^�  t�  ^�      H   ,  v<  `�  v<  a�  w  a�  w  `�  v<  `�      H   ,  v<  ^�  v<  _X  w  _X  w  ^�  v<  ^�      H   ,  s�  `�  s�  a�  t�  a�  t�  `�  s�  `�      H   ,  v<  `   v<  `�  w  `�  w  `   v<  `       H   ,  s�  ^�  s�  _X  t�  _X  t�  ^�  s�  ^�      H   ,  t�  ]�  t�  ^�  ut  ^�  ut  ]�  t�  ]�      H   ,  ut  _X  ut  `   v<  `   v<  _X  ut  _X      H   ,  t�  `�  t�  a�  ut  a�  ut  `�  t�  `�      H   ,  v<  a�  v<  bx  w  bx  w  a�  v<  a�      H   ,  x�  _X  x�  `   y\  `   y\  _X  x�  _X      H   ,  z$  _X  z$  `   z�  `   z�  _X  z$  _X      H   ,  w�  ^�  w�  _X  x�  _X  x�  ^�  w�  ^�      H   ,  }D  bx  }D  c@  ~  c@  ~  bx  }D  bx      H   ,  ||  ^�  ||  _X  }D  _X  }D  ^�  ||  ^�      H   ,  y\  a�  y\  bx  z$  bx  z$  a�  y\  a�      H   ,  ||  bx  ||  c@  }D  c@  }D  bx  ||  bx      H   ,  {�  `   {�  `�  ||  `�  ||  `   {�  `       H   ,  w�  ]   w�  ]�  x�  ]�  x�  ]   w�  ]       H   ,  w�  _X  w�  `   x�  `   x�  _X  w�  _X      H   ,  y\  ^�  y\  _X  z$  _X  z$  ^�  y\  ^�      H   ,  z�  _X  z�  `   {�  `   {�  _X  z�  _X      H   ,  }D  a�  }D  bx  ~  bx  ~  a�  }D  a�      H   ,  x�  ]�  x�  ^�  y\  ^�  y\  ]�  x�  ]�      H   ,  w�  `   w�  `�  x�  `�  x�  `   w�  `       H   ,  }D  `�  }D  a�  ~  a�  ~  `�  }D  `�      H   ,  z�  a�  z�  bx  {�  bx  {�  a�  z�  a�      H   ,  y\  bx  y\  c@  z$  c@  z$  bx  y\  bx      H   ,  {�  _X  {�  `   ||  `   ||  _X  {�  _X      H   ,  x�  `   x�  `�  y\  `�  y\  `   x�  `       H   ,  x�  ^�  x�  _X  y\  _X  y\  ^�  x�  ^�      H   ,  z$  ^�  z$  _X  z�  _X  z�  ^�  z$  ^�      H   ,  ||  _X  ||  `   }D  `   }D  _X  ||  _X      H   ,  x�  bx  x�  c@  y\  c@  y\  bx  x�  bx      H   ,  {�  ]   {�  ]�  ||  ]�  ||  ]   {�  ]       H   ,  }D  `   }D  `�  ~  `�  ~  `   }D  `       H   ,  z$  ]�  z$  ^�  z�  ^�  z�  ]�  z$  ]�      H   ,  z�  ]   z�  ]�  {�  ]�  {�  ]   z�  ]       H   ,  x�  ]   x�  ]�  y\  ]�  y\  ]   x�  ]       H   ,  {�  bx  {�  c@  ||  c@  ||  bx  {�  bx      H   ,  y\  ]�  y\  ^�  z$  ^�  z$  ]�  y\  ]�      H   ,  }D  _X  }D  `   ~  `   ~  _X  }D  _X      H   ,  ||  ]   ||  ]�  }D  ]�  }D  ]   ||  ]       H   ,  x�  a�  x�  bx  y\  bx  y\  a�  x�  a�      H   ,  y\  _X  y\  `   z$  `   z$  _X  y\  _X      H   ,  z�  bx  z�  c@  {�  c@  {�  bx  z�  bx      H   ,  {�  ^�  {�  _X  ||  _X  ||  ^�  {�  ^�      H   ,  z�  ^�  z�  _X  {�  _X  {�  ^�  z�  ^�      H   ,  z$  ]   z$  ]�  z�  ]�  z�  ]   z$  ]       H   ,  }D  ^�  }D  _X  ~  _X  ~  ^�  }D  ^�      H   ,  x�  `�  x�  a�  y\  a�  y\  `�  x�  `�      H   ,  ||  `   ||  `�  }D  `�  }D  `   ||  `       H   ,  w�  a�  w�  bx  x�  bx  x�  a�  w�  a�      H   ,  {�  a�  {�  bx  ||  bx  ||  a�  {�  a�      H   ,  w�  `�  w�  a�  x�  a�  x�  `�  w�  `�      H   ,  w�  ]�  w�  ^�  x�  ^�  x�  ]�  w�  ]�      H   ,  ||  ]�  ||  ^�  }D  ^�  }D  ]�  ||  ]�      H   ,  }D  ]�  }D  ^�  ~  ^�  ~  ]�  }D  ]�      H   ,  z$  `   z$  `�  z�  `�  z�  `   z$  `       H   ,  z$  `�  z$  a�  z�  a�  z�  `�  z$  `�      H   ,  ||  `�  ||  a�  }D  a�  }D  `�  ||  `�      H   ,  w�  bx  w�  c@  x�  c@  x�  bx  w�  bx      H   ,  z$  bx  z$  c@  z�  c@  z�  bx  z$  bx      H   ,  {�  `�  {�  a�  ||  a�  ||  `�  {�  `�      H   ,  y\  `   y\  `�  z$  `�  z$  `   y\  `       H   ,  z�  `�  z�  a�  {�  a�  {�  `�  z�  `�      H   ,  z$  a�  z$  bx  z�  bx  z�  a�  z$  a�      H   ,  z�  `   z�  `�  {�  `�  {�  `   z�  `       H   ,  }D  ]   }D  ]�  ~  ]�  ~  ]   }D  ]       H   ,  y\  ]   y\  ]�  z$  ]�  z$  ]   y\  ]       H   ,  ||  a�  ||  bx  }D  bx  }D  a�  ||  a�      H   ,  z�  ]�  z�  ^�  {�  ^�  {�  ]�  z�  ]�      H   ,  y\  `�  y\  a�  z$  a�  z$  `�  y\  `�      H   ,  {�  ]�  {�  ^�  ||  ^�  ||  ]�  {�  ]�      H   ,  s�  N�  s�  O�  t�  O�  t�  N�  s�  N�      H   ,  ut  N�  ut  O�  v<  O�  v<  N�  ut  N�      H   ,  o�  J@  o�  K  p�  K  p�  J@  o�  J@      H   ,  y\  N�  y\  O�  z$  O�  z$  N�  y\  N�      H   ,  o�  Ix  o�  J@  p�  J@  p�  Ix  o�  Ix      H   ,  rT  N�  rT  O�  s  O�  s  N�  rT  N�      H   ,  o�  K�  o�  L�  p�  L�  p�  K�  o�  K�      H   ,  ||  N�  ||  O�  }D  O�  }D  N�  ||  N�      H   ,  o�  M`  o�  N(  p�  N(  p�  M`  o�  M`      H   ,  q�  N�  q�  O�  rT  O�  rT  N�  q�  N�      H   ,  {�  N�  {�  O�  ||  O�  ||  N�  {�  N�      H   ,  z$  N�  z$  O�  z�  O�  z�  N�  z$  N�      H   ,  o�  K  o�  K�  p�  K�  p�  K  o�  K      H   ,  o�  N(  o�  N�  p�  N�  p�  N(  o�  N(      H   ,  t�  N�  t�  O�  ut  O�  ut  N�  t�  N�      H   ,  w�  N�  w�  O�  x�  O�  x�  N�  w�  N�      H   ,  w  N�  w  O�  w�  O�  w�  N�  w  N�      H   ,  v<  N�  v<  O�  w  O�  w  N�  v<  N�      H   ,  z�  N�  z�  O�  {�  O�  {�  N�  z�  N�      H   ,  }D  N�  }D  O�  ~  O�  ~  N�  }D  N�      H   ,  s  N�  s  O�  s�  O�  s�  N�  s  N�      H   ,  x�  N�  x�  O�  y\  O�  y\  N�  x�  N�      H   ,  o�  L�  o�  M`  p�  M`  p�  L�  o�  L�      H   ,  w  \8  w  ]   w�  ]   w�  \8  w  \8      H   ,  {�  U�  {�  V�  ||  V�  ||  U�  {�  U�      H   ,  w  [p  w  \8  w�  \8  w�  [p  w  [p      H   ,  w  P�  w  QH  w�  QH  w�  P�  w  P�      H   ,  w  Z�  w  [p  w�  [p  w�  Z�  w  Z�      H   ,  w  O�  w  P�  w�  P�  w�  O�  w  O�      H   ,  }D  U�  }D  V�  ~  V�  ~  U�  }D  U�      H   ,  w  Y  w  Y�  w�  Y�  w�  Y  w  Y      H   ,  w  Y�  w  Z�  w�  Z�  w�  Y�  w  Y�      H   ,  ||  U�  ||  V�  }D  V�  }D  U�  ||  U�      H   ,  z$  [p  z$  \8  z�  \8  z�  [p  z$  [p      H   ,  y\  Y�  y\  Z�  z$  Z�  z$  Y�  y\  Y�      H   ,  w�  Z�  w�  [p  x�  [p  x�  Z�  w�  Z�      H   ,  z�  XP  z�  Y  {�  Y  {�  XP  z�  XP      H   ,  z$  Y  z$  Y�  z�  Y�  z�  Y  z$  Y      H   ,  z�  \8  z�  ]   {�  ]   {�  \8  z�  \8      H   ,  y\  \8  y\  ]   z$  ]   z$  \8  y\  \8      H   ,  ||  \8  ||  ]   }D  ]   }D  \8  ||  \8      H   ,  }D  \8  }D  ]   ~  ]   ~  \8  }D  \8      H   ,  w�  Y�  w�  Z�  x�  Z�  x�  Y�  w�  Y�      H   ,  {�  Y  {�  Y�  ||  Y�  ||  Y  {�  Y      H   ,  x�  \8  x�  ]   y\  ]   y\  \8  x�  \8      H   ,  }D  [p  }D  \8  ~  \8  ~  [p  }D  [p      H   ,  ||  [p  ||  \8  }D  \8  }D  [p  ||  [p      H   ,  {�  V�  {�  W�  ||  W�  ||  V�  {�  V�      H   ,  y\  Y  y\  Y�  z$  Y�  z$  Y  y\  Y      H   ,  y\  Z�  y\  [p  z$  [p  z$  Z�  y\  Z�      H   ,  }D  Z�  }D  [p  ~  [p  ~  Z�  }D  Z�      H   ,  x�  [p  x�  \8  y\  \8  y\  [p  x�  [p      H   ,  ||  Z�  ||  [p  }D  [p  }D  Z�  ||  Z�      H   ,  z�  [p  z�  \8  {�  \8  {�  [p  z�  [p      H   ,  w�  Y  w�  Y�  x�  Y�  x�  Y  w�  Y      H   ,  }D  Y�  }D  Z�  ~  Z�  ~  Y�  }D  Y�      H   ,  x�  Z�  x�  [p  y\  [p  y\  Z�  x�  Z�      H   ,  }D  Y  }D  Y�  ~  Y�  ~  Y  }D  Y      H   ,  ||  Y�  ||  Z�  }D  Z�  }D  Y�  ||  Y�      H   ,  z$  XP  z$  Y  z�  Y  z�  XP  z$  XP      H   ,  }D  XP  }D  Y  ~  Y  ~  XP  }D  XP      H   ,  x�  Y�  x�  Z�  y\  Z�  y\  Y�  x�  Y�      H   ,  }D  W�  }D  XP  ~  XP  ~  W�  }D  W�      H   ,  ||  Y  ||  Y�  }D  Y�  }D  Y  ||  Y      H   ,  z�  Z�  z�  [p  {�  [p  {�  Z�  z�  Z�      H   ,  y\  XP  y\  Y  z$  Y  z$  XP  y\  XP      H   ,  }D  V�  }D  W�  ~  W�  ~  V�  }D  V�      H   ,  {�  \8  {�  ]   ||  ]   ||  \8  {�  \8      H   ,  w�  \8  w�  ]   x�  ]   x�  \8  w�  \8      H   ,  {�  XP  {�  Y  ||  Y  ||  XP  {�  XP      H   ,  x�  Y  x�  Y�  y\  Y�  y\  Y  x�  Y      H   ,  ||  XP  ||  Y  }D  Y  }D  XP  ||  XP      H   ,  z�  Y�  z�  Z�  {�  Z�  {�  Y�  z�  Y�      H   ,  x�  XP  x�  Y  y\  Y  y\  XP  x�  XP      H   ,  ||  W�  ||  XP  }D  XP  }D  W�  ||  W�      H   ,  {�  [p  {�  \8  ||  \8  ||  [p  {�  [p      H   ,  {�  Y�  {�  Z�  ||  Z�  ||  Y�  {�  Y�      H   ,  w�  [p  w�  \8  x�  \8  x�  [p  w�  [p      H   ,  ||  V�  ||  W�  }D  W�  }D  V�  ||  V�      H   ,  y\  [p  y\  \8  z$  \8  z$  [p  y\  [p      H   ,  z$  Y�  z$  Z�  z�  Z�  z�  Y�  z$  Y�      H   ,  z$  Z�  z$  [p  z�  [p  z�  Z�  z$  Z�      H   ,  z�  Y  z�  Y�  {�  Y�  {�  Y  z�  Y      H   ,  {�  Z�  {�  [p  ||  [p  ||  Z�  {�  Z�      H   ,  z$  \8  z$  ]   z�  ]   z�  \8  z$  \8      H   ,  {�  W�  {�  XP  ||  XP  ||  W�  {�  W�      H   ,  v<  Y�  v<  Z�  w  Z�  w  Y�  v<  Y�      H   ,  v<  [p  v<  \8  w  \8  w  [p  v<  [p      H   ,  ut  [p  ut  \8  v<  \8  v<  [p  ut  [p      H   ,  v<  \8  v<  ]   w  ]   w  \8  v<  \8      H   ,  t�  [p  t�  \8  ut  \8  ut  [p  t�  [p      H   ,  v<  Z�  v<  [p  w  [p  w  Z�  v<  Z�      H   ,  ut  \8  ut  ]   v<  ]   v<  \8  ut  \8      H   ,  t�  \8  t�  ]   ut  ]   ut  \8  t�  \8      H   ,  ut  Z�  ut  [p  v<  [p  v<  Z�  ut  Z�      H   ,  v<  O�  v<  P�  w  P�  w  O�  v<  O�      H   ,  v<  P�  v<  QH  w  QH  w  P�  v<  P�      H   ,  ut  O�  ut  P�  v<  P�  v<  O�  ut  O�      H   ,  t�  O�  t�  P�  ut  P�  ut  O�  t�  O�      H   ,  s�  O�  s�  P�  t�  P�  t�  O�  s�  O�      H   ,  }D  S�  }D  Th  ~  Th  ~  S�  }D  S�      H   ,  z$  QH  z$  R  z�  R  z�  QH  z$  QH      H   ,  }D  R�  }D  S�  ~  S�  ~  R�  }D  R�      H   ,  ||  Th  ||  U0  }D  U0  }D  Th  ||  Th      H   ,  y\  O�  y\  P�  z$  P�  z$  O�  y\  O�      H   ,  w�  O�  w�  P�  x�  P�  x�  O�  w�  O�      H   ,  }D  R  }D  R�  ~  R�  ~  R  }D  R      H   ,  }D  QH  }D  R  ~  R  ~  QH  }D  QH      H   ,  w�  P�  w�  QH  x�  QH  x�  P�  w�  P�      H   ,  z�  P�  z�  QH  {�  QH  {�  P�  z�  P�      H   ,  {�  O�  {�  P�  ||  P�  ||  O�  {�  O�      H   ,  }D  P�  }D  QH  ~  QH  ~  P�  }D  P�      H   ,  ||  P�  ||  QH  }D  QH  }D  P�  ||  P�      H   ,  }D  O�  }D  P�  ~  P�  ~  O�  }D  O�      H   ,  x�  P�  x�  QH  y\  QH  y\  P�  x�  P�      H   ,  {�  P�  {�  QH  ||  QH  ||  P�  {�  P�      H   ,  }D  U0  }D  U�  ~  U�  ~  U0  }D  U0      H   ,  {�  QH  {�  R  ||  R  ||  QH  {�  QH      H   ,  z$  P�  z$  QH  z�  QH  z�  P�  z$  P�      H   ,  z�  O�  z�  P�  {�  P�  {�  O�  z�  O�      H   ,  z�  QH  z�  R  {�  R  {�  QH  z�  QH      H   ,  x�  O�  x�  P�  y\  P�  y\  O�  x�  O�      H   ,  y\  P�  y\  QH  z$  QH  z$  P�  y\  P�      H   ,  ||  S�  ||  Th  }D  Th  }D  S�  ||  S�      H   ,  }D  Th  }D  U0  ~  U0  ~  Th  }D  Th      H   ,  ||  QH  ||  R  }D  R  }D  QH  ||  QH      H   ,  ||  U0  ||  U�  }D  U�  }D  U0  ||  U0      H   ,  z$  O�  z$  P�  z�  P�  z�  O�  z$  O�      H   ,  ||  O�  ||  P�  }D  P�  }D  O�  ||  O�      H   ,  h�  Ix  h�  J@  i�  J@  i�  Ix  h�  Ix      H   ,  kL  G�  kL  H�  l  H�  l  G�  kL  G�      H   ,  h�  H�  h�  Ix  i�  Ix  i�  H�  h�  H�      H   ,  l�  G�  l�  H�  m�  H�  m�  G�  l�  G�      H   ,  h�  J@  h�  K  i�  K  i�  J@  h�  J@      H   ,  h�  E�  h�  FX  i�  FX  i�  E�  h�  E�      H   ,  h�  FX  h�  G   i�  G   i�  FX  h�  FX      H   ,  j�  G�  j�  H�  kL  H�  kL  G�  j�  G�      H   ,  gd  G�  gd  H�  h,  H�  h,  G�  gd  G�      H   ,  l  G�  l  H�  l�  H�  l�  G�  l  G�      H   ,  e  G�  e  H�  e�  H�  e�  G�  e  G�      H   ,  f�  G�  f�  H�  gd  H�  gd  G�  f�  G�      H   ,  h�  G�  h�  H�  i�  H�  i�  G�  h�  G�      H   ,  h,  G�  h,  H�  h�  H�  h�  G�  h,  G�      H   ,  e�  G�  e�  H�  f�  H�  f�  G�  e�  G�      H   ,  h�  K  h�  K�  i�  K�  i�  K  h�  K      H   ,  h�  G   h�  G�  i�  G�  i�  G   h�  G       H   ,  i�  G�  i�  H�  j�  H�  j�  G�  i�  G�      H   ,  l�  Ix  l�  J@  m�  J@  m�  Ix  l�  Ix      H   ,  nl  H�  nl  Ix  o4  Ix  o4  H�  nl  H�      H   ,  j�  K  j�  K�  kL  K�  kL  K  j�  K      H   ,  kL  H�  kL  Ix  l  Ix  l  H�  kL  H�      H   ,  o4  L�  o4  M`  o�  M`  o�  L�  o4  L�      H   ,  nl  L�  nl  M`  o4  M`  o4  L�  nl  L�      H   ,  l�  L�  l�  M`  m�  M`  m�  L�  l�  L�      H   ,  kL  K�  kL  L�  l  L�  l  K�  kL  K�      H   ,  l�  K�  l�  L�  m�  L�  m�  K�  l�  K�      H   ,  m�  J@  m�  K  nl  K  nl  J@  m�  J@      H   ,  m�  H�  m�  Ix  nl  Ix  nl  H�  m�  H�      H   ,  nl  M`  nl  N(  o4  N(  o4  M`  nl  M`      H   ,  kL  K  kL  K�  l  K�  l  K  kL  K      H   ,  o4  K�  o4  L�  o�  L�  o�  K�  o4  K�      H   ,  j�  J@  j�  K  kL  K  kL  J@  j�  J@      H   ,  nl  Ix  nl  J@  o4  J@  o4  Ix  nl  Ix      H   ,  m�  L�  m�  M`  nl  M`  nl  L�  m�  L�      H   ,  l  K�  l  L�  l�  L�  l�  K�  l  K�      H   ,  kL  J@  kL  K  l  K  l  J@  kL  J@      H   ,  l  L�  l  M`  l�  M`  l�  L�  l  L�      H   ,  j�  K�  j�  L�  kL  L�  kL  K�  j�  K�      H   ,  i�  K  i�  K�  j�  K�  j�  K  i�  K      H   ,  i�  H�  i�  Ix  j�  Ix  j�  H�  i�  H�      H   ,  o4  K  o4  K�  o�  K�  o�  K  o4  K      H   ,  nl  K�  nl  L�  o4  L�  o4  K�  nl  K�      H   ,  l  K  l  K�  l�  K�  l�  K  l  K      H   ,  l  Ix  l  J@  l�  J@  l�  Ix  l  Ix      H   ,  l�  J@  l�  K  m�  K  m�  J@  l�  J@      H   ,  o4  N(  o4  N�  o�  N�  o�  N(  o4  N(      H   ,  m�  K�  m�  L�  nl  L�  nl  K�  m�  K�      H   ,  m�  Ix  m�  J@  nl  J@  nl  Ix  m�  Ix      H   ,  o4  J@  o4  K  o�  K  o�  J@  o4  J@      H   ,  o4  M`  o4  N(  o�  N(  o�  M`  o4  M`      H   ,  l�  H�  l�  Ix  m�  Ix  m�  H�  l�  H�      H   ,  l  H�  l  Ix  l�  Ix  l�  H�  l  H�      H   ,  l�  K  l�  K�  m�  K�  m�  K  l�  K      H   ,  nl  J@  nl  K  o4  K  o4  J@  nl  J@      H   ,  o4  Ix  o4  J@  o�  J@  o�  Ix  o4  Ix      H   ,  i�  J@  i�  K  j�  K  j�  J@  i�  J@      H   ,  m�  K  m�  K�  nl  K�  nl  K  m�  K      H   ,  nl  K  nl  K�  o4  K�  o4  K  nl  K      H   ,  j�  H�  j�  Ix  kL  Ix  kL  H�  j�  H�      H   ,  j�  Ix  j�  J@  kL  J@  kL  Ix  j�  Ix      H   ,  l  J@  l  K  l�  K  l�  J@  l  J@      H   ,  i�  Ix  i�  J@  j�  J@  j�  Ix  i�  Ix      H   ,  m�  M`  m�  N(  nl  N(  nl  M`  m�  M`      H   ,  kL  Ix  kL  J@  l  J@  l  Ix  kL  Ix      H   ,  f�  H�  f�  Ix  gd  Ix  gd  H�  f�  H�      H   ,  h,  Ix  h,  J@  h�  J@  h�  Ix  h,  Ix      H   ,  e�  H�  e�  Ix  f�  Ix  f�  H�  e�  H�      H   ,  f�  Ix  f�  J@  gd  J@  gd  Ix  f�  Ix      H   ,  h,  H�  h,  Ix  h�  Ix  h�  H�  h,  H�      H   ,  gd  J@  gd  K  h,  K  h,  J@  gd  J@      H   ,  h,  J@  h,  K  h�  K  h�  J@  h,  J@      H   ,  gd  H�  gd  Ix  h,  Ix  h,  H�  gd  H�      H   ,  gd  Ix  gd  J@  h,  J@  h,  Ix  gd  Ix      H   ,  e�  D   e�  D�  f�  D�  f�  D   e�  D       H   ,  dD  A�  dD  Bp  e  Bp  e  A�  dD  A�      H   ,  f�  Bp  f�  C8  gd  C8  gd  Bp  f�  Bp      H   ,  f�  C8  f�  D   gd  D   gd  C8  f�  C8      H   ,  e  C8  e  D   e�  D   e�  C8  e  C8      H   ,  dD  G   dD  G�  e  G�  e  G   dD  G       H   ,  dD  C8  dD  D   e  D   e  C8  dD  C8      H   ,  c|  C8  c|  D   dD  D   dD  C8  c|  C8      H   ,  b�  D   b�  D�  c|  D�  c|  D   b�  D       H   ,  gd  D   gd  D�  h,  D�  h,  D   gd  D       H   ,  f�  G   f�  G�  gd  G�  gd  G   f�  G       H   ,  e�  A�  e�  Bp  f�  Bp  f�  A�  e�  A�      H   ,  c|  D�  c|  E�  dD  E�  dD  D�  c|  D�      H   ,  h,  G   h,  G�  h�  G�  h�  G   h,  G       H   ,  e  G   e  G�  e�  G�  e�  G   e  G       H   ,  dD  Bp  dD  C8  e  C8  e  Bp  dD  Bp      H   ,  gd  E�  gd  FX  h,  FX  h,  E�  gd  E�      H   ,  gd  G   gd  G�  h,  G�  h,  G   gd  G       H   ,  h,  FX  h,  G   h�  G   h�  FX  h,  FX      H   ,  e�  E�  e�  FX  f�  FX  f�  E�  e�  E�      H   ,  b�  C8  b�  D   c|  D   c|  C8  b�  C8      H   ,  dD  D�  dD  E�  e  E�  e  D�  dD  D�      H   ,  h,  E�  h,  FX  h�  FX  h�  E�  h,  E�      H   ,  c|  FX  c|  G   dD  G   dD  FX  c|  FX      H   ,  e  A�  e  Bp  e�  Bp  e�  A�  e  A�      H   ,  c|  Bp  c|  C8  dD  C8  dD  Bp  c|  Bp      H   ,  h,  D�  h,  E�  h�  E�  h�  D�  h,  D�      H   ,  f�  FX  f�  G   gd  G   gd  FX  f�  FX      H   ,  e�  Bp  e�  C8  f�  C8  f�  Bp  e�  Bp      H   ,  f�  D   f�  D�  gd  D�  gd  D   f�  D       H   ,  e�  G   e�  G�  f�  G�  f�  G   e�  G       H   ,  e  D   e  D�  e�  D�  e�  D   e  D       H   ,  e  FX  e  G   e�  G   e�  FX  e  FX      H   ,  dD  FX  dD  G   e  G   e  FX  dD  FX      H   ,  e�  C8  e�  D   f�  D   f�  C8  e�  C8      H   ,  b�  Bp  b�  C8  c|  C8  c|  Bp  b�  Bp      H   ,  b�  A�  b�  Bp  c|  Bp  c|  A�  b�  A�      H   ,  gd  D�  gd  E�  h,  E�  h,  D�  gd  D�      H   ,  f�  E�  f�  FX  gd  FX  gd  E�  f�  E�      H   ,  b�  D�  b�  E�  c|  E�  c|  D�  b�  D�      H   ,  c|  E�  c|  FX  dD  FX  dD  E�  c|  E�      H   ,  gd  FX  gd  G   h,  G   h,  FX  gd  FX      H   ,  c|  A�  c|  Bp  dD  Bp  dD  A�  c|  A�      H   ,  dD  D   dD  D�  e  D�  e  D   dD  D       H   ,  e�  FX  e�  G   f�  G   f�  FX  e�  FX      H   ,  e�  D�  e�  E�  f�  E�  f�  D�  e�  D�      H   ,  e  E�  e  FX  e�  FX  e�  E�  e  E�      H   ,  c|  D   c|  D�  dD  D�  dD  D   c|  D       H   ,  dD  E�  dD  FX  e  FX  e  E�  dD  E�      H   ,  e  D�  e  E�  e�  E�  e�  D�  e  D�      H   ,  f�  D�  f�  E�  gd  E�  gd  D�  f�  D�      H   ,  e  Bp  e  C8  e�  C8  e�  Bp  e  Bp      H   ,  j�  G   j�  G�  kL  G�  kL  G   j�  G       H   ,  i�  FX  i�  G   j�  G   j�  FX  i�  FX      H   ,  j�  FX  j�  G   kL  G   kL  FX  j�  FX      H   ,  i�  G   i�  G�  j�  G�  j�  G   i�  G       H   ,  kL  G   kL  G�  l  G�  l  G   kL  G       H   ,  s�  K  s�  K�  t�  K�  t�  K  s�  K      H   ,  {�  M`  {�  N(  ||  N(  ||  M`  {�  M`      H   ,  s�  M`  s�  N(  t�  N(  t�  M`  s�  M`      H   ,  q�  K�  q�  L�  rT  L�  rT  K�  q�  K�      H   ,  y\  N(  y\  N�  z$  N�  z$  N(  y\  N(      H   ,  t�  K  t�  K�  ut  K�  ut  K  t�  K      H   ,  p�  J@  p�  K  q�  K  q�  J@  p�  J@      H   ,  w  M`  w  N(  w�  N(  w�  M`  w  M`      H   ,  q�  N(  q�  N�  rT  N�  rT  N(  q�  N(      H   ,  z$  L�  z$  M`  z�  M`  z�  L�  z$  L�      H   ,  x�  M`  x�  N(  y\  N(  y\  M`  x�  M`      H   ,  p�  K  p�  K�  q�  K�  q�  K  p�  K      H   ,  v<  L�  v<  M`  w  M`  w  L�  v<  L�      H   ,  p�  N(  p�  N�  q�  N�  q�  N(  p�  N(      H   ,  rT  K  rT  K�  s  K�  s  K  rT  K      H   ,  v<  M`  v<  N(  w  N(  w  M`  v<  M`      H   ,  z�  N(  z�  N�  {�  N�  {�  N(  z�  N(      H   ,  w�  M`  w�  N(  x�  N(  x�  M`  w�  M`      H   ,  ut  M`  ut  N(  v<  N(  v<  M`  ut  M`      H   ,  s  K  s  K�  s�  K�  s�  K  s  K      H   ,  w  K�  w  L�  w�  L�  w�  K�  w  K�      H   ,  s�  K�  s�  L�  t�  L�  t�  K�  s�  K�      H   ,  rT  M`  rT  N(  s  N(  s  M`  rT  M`      H   ,  q�  M`  q�  N(  rT  N(  rT  M`  q�  M`      H   ,  ||  N(  ||  N�  }D  N�  }D  N(  ||  N(      H   ,  q�  K  q�  K�  rT  K�  rT  K  q�  K      H   ,  p�  M`  p�  N(  q�  N(  q�  M`  p�  M`      H   ,  rT  J@  rT  K  s  K  s  J@  rT  J@      H   ,  z$  N(  z$  N�  z�  N�  z�  N(  z$  N(      H   ,  y\  M`  y\  N(  z$  N(  z$  M`  y\  M`      H   ,  s  N(  s  N�  s�  N�  s�  N(  s  N(      H   ,  }D  N(  }D  N�  ~  N�  ~  N(  }D  N(      H   ,  s  M`  s  N(  s�  N(  s�  M`  s  M`      H   ,  {�  N(  {�  N�  ||  N�  ||  N(  {�  N(      H   ,  w  L�  w  M`  w�  M`  w�  L�  w  L�      H   ,  w  N(  w  N�  w�  N�  w�  N(  w  N(      H   ,  }D  M`  }D  N(  ~  N(  ~  M`  }D  M`      H   ,  z�  M`  z�  N(  {�  N(  {�  M`  z�  M`      H   ,  v<  N(  v<  N�  w  N�  w  N(  v<  N(      H   ,  p�  K�  p�  L�  q�  L�  q�  K�  p�  K�      H   ,  y\  L�  y\  M`  z$  M`  z$  L�  y\  L�      H   ,  w�  L�  w�  M`  x�  M`  x�  L�  w�  L�      H   ,  t�  N(  t�  N�  ut  N�  ut  N(  t�  N(      H   ,  rT  L�  rT  M`  s  M`  s  L�  rT  L�      H   ,  ut  N(  ut  N�  v<  N�  v<  N(  ut  N(      H   ,  ||  M`  ||  N(  }D  N(  }D  M`  ||  M`      H   ,  q�  L�  q�  M`  rT  M`  rT  L�  q�  L�      H   ,  t�  M`  t�  N(  ut  N(  ut  M`  t�  M`      H   ,  s�  L�  s�  M`  t�  M`  t�  L�  s�  L�      H   ,  ut  L�  ut  M`  v<  M`  v<  L�  ut  L�      H   ,  z$  M`  z$  N(  z�  N(  z�  M`  z$  M`      H   ,  p�  L�  p�  M`  q�  M`  q�  L�  p�  L�      H   ,  s�  N(  s�  N�  t�  N�  t�  N(  s�  N(      H   ,  t�  L�  t�  M`  ut  M`  ut  L�  t�  L�      H   ,  w�  K�  w�  L�  x�  L�  x�  K�  w�  K�      H   ,  q�  J@  q�  K  rT  K  rT  J@  q�  J@      H   ,  s  K�  s  L�  s�  L�  s�  K�  s  K�      H   ,  x�  N(  x�  N�  y\  N�  y\  N(  x�  N(      H   ,  ut  K�  ut  L�  v<  L�  v<  K�  ut  K�      H   ,  v<  K�  v<  L�  w  L�  w  K�  v<  K�      H   ,  w�  N(  w�  N�  x�  N�  x�  N(  w�  N(      H   ,  x�  L�  x�  M`  y\  M`  y\  L�  x�  L�      H   ,  rT  K�  rT  L�  s  L�  s  K�  rT  K�      H   ,  rT  N(  rT  N�  s  N�  s  N(  rT  N(      H   ,  t�  K�  t�  L�  ut  L�  ut  K�  t�  K�      H   ,  s  L�  s  M`  s�  M`  s�  L�  s  L�      H   ,  ��  N�  ��  O�  �L  O�  �L  N�  ��  N�      H   ,  �<  N�  �<  O�  �  O�  �  N�  �<  N�      H   ,  �T  G   �T  G�  �  G�  �  G   �T  G       H   ,  �\  N�  �\  O�  �$  O�  �$  N�  �\  N�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �T  FX  �T  G   �  G   �  FX  �T  FX      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �T  E�  �T  FX  �  FX  �  E�  �T  E�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �T  D�  �T  E�  �  E�  �  D�  �T  D�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  ��  N�  ��  O�  �t  O�  �t  N�  ��  N�      H   ,  �  N�  �  O�  ��  O�  ��  N�  �  N�      H   ,  �T  D   �T  D�  �  D�  �  D   �T  D       H   ,  �,  N�  �,  O�  ��  O�  ��  N�  �,  N�      H   ,  �L  N�  �L  O�  �  O�  �  N�  �L  N�      H   ,  �T  C8  �T  D   �  D   �  C8  �T  C8      H   ,  �T  Bp  �T  C8  �  C8  �  Bp  �T  Bp      H   ,  �T  A�  �T  Bp  �  Bp  �  A�  �T  A�      H   ,  ��  N�  ��  O�  �l  O�  �l  N�  ��  N�      H   ,  �T  S�  �T  Th  �  Th  �  S�  �T  S�      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �T  R�  �T  S�  �  S�  �  R�  �T  R�      H   ,  �t  N�  �t  O�  �<  O�  �<  N�  �t  N�      H   ,  �T  R  �T  R�  �  R�  �  R  �T  R      H   ,  ��  N�  ��  O�  ��  O�  ��  N�  ��  N�      H   ,  �T  QH  �T  R  �  R  �  QH  �T  QH      H   ,  �4  N�  �4  O�  ��  O�  ��  N�  �4  N�      H   ,  �T  P�  �T  QH  �  QH  �  P�  �T  P�      H   ,  ��  N�  ��  O�  �\  O�  �\  N�  ��  N�      H   ,  ~�  N�  ~�  O�  �  O�  �  N�  ~�  N�      H   ,  �T  O�  �T  P�  �  P�  �  O�  �T  O�      H   ,  �  N�  �  O�  �d  O�  �d  N�  �  N�      H   ,  �T  J@  �T  K  �  K  �  J@  �T  J@      H   ,  �  N�  �  O�  ��  O�  ��  N�  �  N�      H   ,  �T  Ix  �T  J@  �  J@  �  Ix  �T  Ix      H   ,  �T  H�  �T  Ix  �  Ix  �  H�  �T  H�      H   ,  �T  G�  �T  H�  �  H�  �  G�  �T  G�      H   ,  ~  N�  ~  O�  ~�  O�  ~�  N�  ~  N�      H   ,  �d  N�  �d  O�  �,  O�  �,  N�  �d  N�      H   ,  �l  N�  �l  O�  �4  O�  �4  N�  �l  N�      H   ,  �\  O�  �\  P�  �$  P�  �$  O�  �\  O�      H   ,  �$  U�  �$  V�  ��  V�  ��  U�  �$  U�      H   ,  ��  U�  ��  V�  �|  V�  �|  U�  ��  U�      H   ,  �\  W�  �\  XP  �$  XP  �$  W�  �\  W�      H   ,  �\  V�  �\  W�  �$  W�  �$  V�  �\  V�      H   ,  ��  U�  ��  V�  ��  V�  ��  U�  ��  U�      H   ,  �\  U�  �\  V�  �$  V�  �$  U�  �\  U�      H   ,  �|  U�  �|  V�  �D  V�  �D  U�  �|  U�      H   ,  �\  P�  �\  QH  �$  QH  �$  P�  �\  P�      H   ,  �\  U0  �\  U�  �$  U�  �$  U0  �\  U0      H   ,  �D  U�  �D  V�  �  V�  �  U�  �D  U�      H   ,  �\  Th  �\  U0  �$  U0  �$  Th  �\  Th      H   ,  �\  S�  �\  Th  �$  Th  �$  S�  �\  S�      H   ,  �\  R�  �\  S�  �$  S�  �$  R�  �\  R�      H   ,  ��  U�  ��  V�  �\  V�  �\  U�  ��  U�      H   ,  �\  R  �\  R�  �$  R�  �$  R  �\  R      H   ,  �\  QH  �\  R  �$  R  �$  QH  �\  QH      H   ,  �D  \8  �D  ]   �  ]   �  \8  �D  \8      H   ,  ��  W�  ��  XP  ��  XP  ��  W�  ��  W�      H   ,  �  Y  �  Y�  ��  Y�  ��  Y  �  Y      H   ,  ��  Y  ��  Y�  �d  Y�  �d  Y  ��  Y      H   ,  ��  XP  ��  Y  ��  Y  ��  XP  ��  XP      H   ,  �D  [p  �D  \8  �  \8  �  [p  �D  [p      H   ,  �|  [p  �|  \8  �D  \8  �D  [p  �|  [p      H   ,  ��  \8  ��  ]   �d  ]   �d  \8  ��  \8      H   ,  �D  Z�  �D  [p  �  [p  �  Z�  �D  Z�      H   ,  �  Z�  �  [p  ��  [p  ��  Z�  �  Z�      H   ,  ��  Y�  ��  Z�  ��  Z�  ��  Y�  ��  Y�      H   ,  �D  Y�  �D  Z�  �  Z�  �  Y�  �D  Y�      H   ,  �|  V�  �|  W�  �D  W�  �D  V�  �|  V�      H   ,  ��  Y�  ��  Z�  ��  Z�  ��  Y�  ��  Y�      H   ,  �D  Y  �D  Y�  �  Y�  �  Y  �D  Y      H   ,  �|  Z�  �|  [p  �D  [p  �D  Z�  �|  Z�      H   ,  �  XP  �  Y  ��  Y  ��  XP  �  XP      H   ,  ��  W�  ��  XP  �|  XP  �|  W�  ��  W�      H   ,  �D  XP  �D  Y  �  Y  �  XP  �D  XP      H   ,  ��  Y�  ��  Z�  �|  Z�  �|  Y�  ��  Y�      H   ,  �|  XP  �|  Y  �D  Y  �D  XP  �|  XP      H   ,  �D  W�  �D  XP  �  XP  �  W�  �D  W�      H   ,  �  W�  �  XP  ��  XP  ��  W�  �  W�      H   ,  �$  V�  �$  W�  ��  W�  ��  V�  �$  V�      H   ,  ��  [p  ��  \8  �d  \8  �d  [p  ��  [p      H   ,  �D  V�  �D  W�  �  W�  �  V�  �D  V�      H   ,  �|  Y  �|  Y�  �D  Y�  �D  Y  �|  Y      H   ,  ��  \8  ��  ]   ��  ]   ��  \8  ��  \8      H   ,  ��  [p  ��  \8  �|  \8  �|  [p  ��  [p      H   ,  ��  XP  ��  Y  ��  Y  ��  XP  ��  XP      H   ,  �|  W�  �|  XP  �D  XP  �D  W�  �|  W�      H   ,  ��  Y  ��  Y�  ��  Y�  ��  Y  ��  Y      H   ,  �  Y�  �  Z�  ��  Z�  ��  Y�  �  Y�      H   ,  ��  Y  ��  Y�  ��  Y�  ��  Y  ��  Y      H   ,  �|  \8  �|  ]   �D  ]   �D  \8  �|  \8      H   ,  ��  Y  ��  Y�  �|  Y�  �|  Y  ��  Y      H   ,  ��  Z�  ��  [p  �d  [p  �d  Z�  ��  Z�      H   ,  ��  [p  ��  \8  ��  \8  ��  [p  ��  [p      H   ,  ��  Z�  ��  [p  �|  [p  �|  Z�  ��  Z�      H   ,  ��  Y�  ��  Z�  �d  Z�  �d  Y�  ��  Y�      H   ,  ��  W�  ��  XP  ��  XP  ��  W�  ��  W�      H   ,  �|  Y�  �|  Z�  �D  Z�  �D  Y�  �|  Y�      H   ,  �$  Y  �$  Y�  ��  Y�  ��  Y  �$  Y      H   ,  �$  W�  �$  XP  ��  XP  ��  W�  �$  W�      H   ,  �  \8  �  ]   ��  ]   ��  \8  �  \8      H   ,  ��  V�  ��  W�  ��  W�  ��  V�  ��  V�      H   ,  �  V�  �  W�  ��  W�  ��  V�  �  V�      H   ,  ��  V�  ��  W�  �|  W�  �|  V�  ��  V�      H   ,  �  [p  �  \8  ��  \8  ��  [p  �  [p      H   ,  ��  Z�  ��  [p  ��  [p  ��  Z�  ��  Z�      H   ,  ��  XP  ��  Y  �|  Y  �|  XP  ��  XP      H   ,  �$  XP  �$  Y  ��  Y  ��  XP  �$  XP      H   ,  �  R�  �  S�  ��  S�  ��  R�  �  R�      H   ,  �  R  �  R�  ��  R�  ��  R  �  R      H   ,  ��  R  ��  R�  �t  R�  �t  R  ��  R      H   ,  ��  Th  ��  U0  ��  U0  ��  Th  ��  Th      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  �  R  �  R�  ��  R�  ��  R  �  R      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �  QH  �  R  ��  R  ��  QH  �  QH      H   ,  �t  QH  �t  R  �<  R  �<  QH  �t  QH      H   ,  �  O�  �  P�  ��  P�  ��  O�  �  O�      H   ,  ��  R�  ��  S�  �t  S�  �t  R�  ��  R�      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  �  P�  �  QH  ��  QH  ��  P�  �  P�      H   ,  �  S�  �  Th  ��  Th  ��  S�  �  S�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �  O�  �  P�  ��  P�  ��  O�  �  O�      H   ,  ��  O�  ��  P�  �t  P�  �t  O�  ��  O�      H   ,  ��  R�  ��  S�  �\  S�  �\  R�  ��  R�      H   ,  �<  S�  �<  Th  �  Th  �  S�  �<  S�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ��  Th  ��  U0  �\  U0  �\  Th  ��  Th      H   ,  ��  P�  ��  QH  �\  QH  �\  P�  ��  P�      H   ,  �t  R  �t  R�  �<  R�  �<  R  �t  R      H   ,  ��  QH  ��  R  �t  R  �t  QH  ��  QH      H   ,  �<  R�  �<  S�  �  S�  �  R�  �<  R�      H   ,  �t  P�  �t  QH  �<  QH  �<  P�  �t  P�      H   ,  �t  S�  �t  Th  �<  Th  �<  S�  �t  S�      H   ,  �  QH  �  R  ��  R  ��  QH  �  QH      H   ,  �<  R  �<  R�  �  R�  �  R  �<  R      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  U0  ��  U�  �\  U�  �\  U0  ��  U0      H   ,  �<  QH  �<  R  �  R  �  QH  �<  QH      H   ,  �  R�  �  S�  ��  S�  ��  R�  �  R�      H   ,  ��  S�  ��  Th  �\  Th  �\  S�  ��  S�      H   ,  ��  O�  ��  P�  �\  P�  �\  O�  ��  O�      H   ,  �<  P�  �<  QH  �  QH  �  P�  �<  P�      H   ,  ��  R  ��  R�  �\  R�  �\  R  ��  R      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  �t  R�  �t  S�  �<  S�  �<  R�  �t  R�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  �t  O�  �t  P�  �<  P�  �<  O�  �t  O�      H   ,  �  S�  �  Th  ��  Th  ��  S�  �  S�      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �  P�  �  QH  ��  QH  ��  P�  �  P�      H   ,  �<  O�  �<  P�  �  P�  �  O�  �<  O�      H   ,  ��  P�  ��  QH  �t  QH  �t  P�  ��  P�      H   ,  ��  S�  ��  Th  �t  Th  �t  S�  ��  S�      H   ,  ��  QH  ��  R  �\  R  �\  QH  ��  QH      H   ,  ��  U0  ��  U�  �|  U�  �|  U0  ��  U0      H   ,  ��  P�  ��  QH  �|  QH  �|  P�  ��  P�      H   ,  ��  Th  ��  U0  �|  U0  �|  Th  ��  Th      H   ,  ��  Th  ��  U0  �d  U0  �d  Th  ��  Th      H   ,  �  P�  �  QH  ��  QH  ��  P�  �  P�      H   ,  �$  Th  �$  U0  ��  U0  ��  Th  �$  Th      H   ,  �|  R  �|  R�  �D  R�  �D  R  �|  R      H   ,  �D  Th  �D  U0  �  U0  �  Th  �D  Th      H   ,  �  R�  �  S�  ��  S�  ��  R�  �  R�      H   ,  �$  R�  �$  S�  ��  S�  ��  R�  �$  R�      H   ,  ��  P�  ��  QH  �d  QH  �d  P�  ��  P�      H   ,  ��  R�  ��  S�  �|  S�  �|  R�  ��  R�      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �$  P�  �$  QH  ��  QH  ��  P�  �$  P�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  �|  Th  �|  U0  �D  U0  �D  Th  �|  Th      H   ,  �  QH  �  R  ��  R  ��  QH  �  QH      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  �D  S�  �D  Th  �  Th  �  S�  �D  S�      H   ,  ��  R  ��  R�  �|  R�  �|  R  ��  R      H   ,  ��  R  ��  R�  �d  R�  �d  R  ��  R      H   ,  ��  Th  ��  U0  ��  U0  ��  Th  ��  Th      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  �|  R�  �|  S�  �D  S�  �D  R�  �|  R�      H   ,  �D  R�  �D  S�  �  S�  �  R�  �D  R�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  U0  ��  U�  ��  U�  ��  U0  ��  U0      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  �D  R  �D  R�  �  R�  �  R  �D  R      H   ,  �|  S�  �|  Th  �D  Th  �D  S�  �|  S�      H   ,  ��  QH  ��  R  �|  R  �|  QH  ��  QH      H   ,  ��  S�  ��  Th  �d  Th  �d  S�  ��  S�      H   ,  �D  QH  �D  R  �  R  �  QH  �D  QH      H   ,  ��  Th  ��  U0  ��  U0  ��  Th  ��  Th      H   ,  ��  S�  ��  Th  �|  Th  �|  S�  ��  S�      H   ,  �$  S�  �$  Th  ��  Th  ��  S�  �$  S�      H   ,  �|  QH  �|  R  �D  R  �D  QH  �|  QH      H   ,  �|  P�  �|  QH  �D  QH  �D  P�  �|  P�      H   ,  �  S�  �  Th  ��  Th  ��  S�  �  S�      H   ,  �  R  �  R�  ��  R�  ��  R  �  R      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �D  P�  �D  QH  �  QH  �  P�  �D  P�      H   ,  ��  QH  ��  R  �d  R  �d  QH  ��  QH      H   ,  ��  O�  ��  P�  �|  P�  �|  O�  ��  O�      H   ,  �|  U0  �|  U�  �D  U�  �D  U0  �|  U0      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  �$  R  �$  R�  ��  R�  ��  R  �$  R      H   ,  �|  O�  �|  P�  �D  P�  �D  O�  �|  O�      H   ,  �$  QH  �$  R  ��  R  ��  QH  �$  QH      H   ,  �$  O�  �$  P�  ��  P�  ��  O�  �$  O�      H   ,  �$  U0  �$  U�  ��  U�  ��  U0  �$  U0      H   ,  ��  R�  ��  S�  �d  S�  �d  R�  ��  R�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �D  U0  �D  U�  �  U�  �  U0  �D  U0      H   ,  �  Th  �  U0  ��  U0  ��  Th  �  Th      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �d  U�  �d  V�  �,  V�  �,  U�  �d  U�      H   ,  �L  P�  �L  QH  �  QH  �  P�  �L  P�      H   ,  �  U�  �  V�  �d  V�  �d  U�  �  U�      H   ,  �L  O�  �L  P�  �  P�  �  O�  �L  O�      H   ,  �L  R�  �L  S�  �  S�  �  R�  �L  R�      H   ,  ~�  U�  ~�  V�  �  V�  �  U�  ~�  U�      H   ,  ~  U�  ~  V�  ~�  V�  ~�  U�  ~  U�      H   ,  �L  R  �L  R�  �  R�  �  R  �L  R      H   ,  �L  QH  �L  R  �  R  �  QH  �L  QH      H   ,  ~  Z�  ~  [p  ~�  [p  ~�  Z�  ~  Z�      H   ,  �d  \8  �d  ]   �,  ]   �,  \8  �d  \8      H   ,  ~�  XP  ~�  Y  �  Y  �  XP  ~�  XP      H   ,  �,  [p  �,  \8  ��  \8  ��  [p  �,  [p      H   ,  �  W�  �  XP  �d  XP  �d  W�  �  W�      H   ,  ~  \8  ~  ]   ~�  ]   ~�  \8  ~  \8      H   ,  �  V�  �  W�  �d  W�  �d  V�  �  V�      H   ,  ~�  Z�  ~�  [p  �  [p  �  Z�  ~�  Z�      H   ,  ~  W�  ~  XP  ~�  XP  ~�  W�  ~  W�      H   ,  �d  [p  �d  \8  �,  \8  �,  [p  �d  [p      H   ,  ~�  Y  ~�  Y�  �  Y�  �  Y  ~�  Y      H   ,  �,  \8  �,  ]   ��  ]   ��  \8  �,  \8      H   ,  ~  Y  ~  Y�  ~�  Y�  ~�  Y  ~  Y      H   ,  �  Z�  �  [p  �d  [p  �d  Z�  �  Z�      H   ,  ~  Y�  ~  Z�  ~�  Z�  ~�  Y�  ~  Y�      H   ,  �  [p  �  \8  �d  \8  �d  [p  �  [p      H   ,  �  Y�  �  Z�  �d  Z�  �d  Y�  �  Y�      H   ,  ~�  V�  ~�  W�  �  W�  �  V�  ~�  V�      H   ,  ~�  W�  ~�  XP  �  XP  �  W�  ~�  W�      H   ,  �  XP  �  Y  �d  Y  �d  XP  �  XP      H   ,  ~�  Y�  ~�  Z�  �  Z�  �  Y�  ~�  Y�      H   ,  ~  XP  ~  Y  ~�  Y  ~�  XP  ~  XP      H   ,  ~  V�  ~  W�  ~�  W�  ~�  V�  ~  V�      H   ,  ~�  [p  ~�  \8  �  \8  �  [p  ~�  [p      H   ,  �d  Z�  �d  [p  �,  [p  �,  Z�  �d  Z�      H   ,  ~�  \8  ~�  ]   �  ]   �  \8  ~�  \8      H   ,  ~  [p  ~  \8  ~�  \8  ~�  [p  ~  [p      H   ,  �  \8  �  ]   �d  ]   �d  \8  �  \8      H   ,  ~  S�  ~  Th  ~�  Th  ~�  S�  ~  S�      H   ,  �d  S�  �d  Th  �,  Th  �,  S�  �d  S�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  �,  P�  �,  QH  ��  QH  ��  P�  �,  P�      H   ,  ~  Th  ~  U0  ~�  U0  ~�  Th  ~  Th      H   ,  �d  Th  �d  U0  �,  U0  �,  Th  �d  Th      H   ,  ~�  S�  ~�  Th  �  Th  �  S�  ~�  S�      H   ,  �d  R  �d  R�  �,  R�  �,  R  �d  R      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ~  U0  ~  U�  ~�  U�  ~�  U0  ~  U0      H   ,  ~  R�  ~  S�  ~�  S�  ~�  R�  ~  R�      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  �  QH  �  R  �d  R  �d  QH  �  QH      H   ,  ��  QH  ��  R  �L  R  �L  QH  ��  QH      H   ,  ~�  R  ~�  R�  �  R�  �  R  ~�  R      H   ,  �,  R�  �,  S�  ��  S�  ��  R�  �,  R�      H   ,  �  R�  �  S�  �d  S�  �d  R�  �  R�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ~  O�  ~  P�  ~�  P�  ~�  O�  ~  O�      H   ,  �d  O�  �d  P�  �,  P�  �,  O�  �d  O�      H   ,  �,  O�  �,  P�  ��  P�  ��  O�  �,  O�      H   ,  ~�  U0  ~�  U�  �  U�  �  U0  ~�  U0      H   ,  �d  R�  �d  S�  �,  S�  �,  R�  �d  R�      H   ,  ~�  P�  ~�  QH  �  QH  �  P�  ~�  P�      H   ,  �  P�  �  QH  �d  QH  �d  P�  �  P�      H   ,  ~�  Th  ~�  U0  �  U0  �  Th  ~�  Th      H   ,  �,  QH  �,  R  ��  R  ��  QH  �,  QH      H   ,  �d  P�  �d  QH  �,  QH  �,  P�  �d  P�      H   ,  �  O�  �  P�  �d  P�  �d  O�  �  O�      H   ,  ~�  QH  ~�  R  �  R  �  QH  ~�  QH      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  �,  S�  �,  Th  ��  Th  ��  S�  �,  S�      H   ,  �  U0  �  U�  �d  U�  �d  U0  �  U0      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �d  QH  �d  R  �,  R  �,  QH  �d  QH      H   ,  ��  R  ��  R�  �L  R�  �L  R  ��  R      H   ,  ~  R  ~  R�  ~�  R�  ~�  R  ~  R      H   ,  ~�  R�  ~�  S�  �  S�  �  R�  ~�  R�      H   ,  ��  R�  ��  S�  �L  S�  �L  R�  ��  R�      H   ,  ��  O�  ��  P�  �L  P�  �L  O�  ��  O�      H   ,  �  R  �  R�  �d  R�  �d  R  �  R      H   ,  ��  P�  ��  QH  �L  QH  �L  P�  ��  P�      H   ,  �  Th  �  U0  �d  U0  �d  Th  �  Th      H   ,  �d  U0  �d  U�  �,  U�  �,  U0  �d  U0      H   ,  �,  R  �,  R�  ��  R�  ��  R  �,  R      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  ~�  O�  ~�  P�  �  P�  �  O�  ~�  O�      H   ,  ~  P�  ~  QH  ~�  QH  ~�  P�  ~  P�      H   ,  �  S�  �  Th  �d  Th  �d  S�  �  S�      H   ,  ~  QH  ~  R  ~�  R  ~�  QH  ~  QH      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  ��  QH  ��  R  �T  R  �T  QH  ��  QH      H   ,  �l  R  �l  R�  �4  R�  �4  R  �l  R      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ��  P�  ��  QH  �l  QH  �l  P�  ��  P�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  R�  ��  S�  �T  S�  �T  R�  ��  R�      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  O�  ��  P�  ��  P�  ��  O�  ��  O�      H   ,  �4  R  �4  R�  ��  R�  ��  R  �4  R      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �  O�  �  P�  ��  P�  ��  O�  �  O�      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �l  QH  �l  R  �4  R  �4  QH  �l  QH      H   ,  �4  R�  �4  S�  ��  S�  ��  R�  �4  R�      H   ,  ��  QH  ��  R  �l  R  �l  QH  ��  QH      H   ,  ��  R�  ��  S�  �l  S�  �l  R�  ��  R�      H   ,  �4  O�  �4  P�  ��  P�  ��  O�  �4  O�      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  �l  S�  �l  Th  �4  Th  �4  S�  �l  S�      H   ,  ��  R  ��  R�  ��  R�  ��  R  ��  R      H   ,  �4  P�  �4  QH  ��  QH  ��  P�  �4  P�      H   ,  �  R�  �  S�  ��  S�  ��  R�  �  R�      H   ,  ��  R  ��  R�  �l  R�  �l  R  ��  R      H   ,  �l  R�  �l  S�  �4  S�  �4  R�  �l  R�      H   ,  �  QH  �  R  ��  R  ��  QH  �  QH      H   ,  ��  R�  ��  S�  ��  S�  ��  R�  ��  R�      H   ,  ��  O�  ��  P�  �T  P�  �T  O�  ��  O�      H   ,  ��  S�  ��  Th  ��  Th  ��  S�  ��  S�      H   ,  ��  R  ��  R�  �T  R�  �T  R  ��  R      H   ,  �4  S�  �4  Th  ��  Th  ��  S�  �4  S�      H   ,  �  P�  �  QH  ��  QH  ��  P�  �  P�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  �  R  �  R�  ��  R�  ��  R  �  R      H   ,  �l  P�  �l  QH  �4  QH  �4  P�  �l  P�      H   ,  ��  P�  ��  QH  ��  QH  ��  P�  ��  P�      H   ,  ��  P�  ��  QH  �T  QH  �T  P�  ��  P�      H   ,  ��  O�  ��  P�  �l  P�  �l  O�  ��  O�      H   ,  �4  QH  �4  R  ��  R  ��  QH  �4  QH      H   ,  �l  O�  �l  P�  �4  P�  �4  O�  �l  O�      H   ,  ��  QH  ��  R  ��  R  ��  QH  ��  QH      H   ,  ��  S�  ��  Th  �T  Th  �T  S�  ��  S�      H   ,  �L  H�  �L  Ix  �  Ix  �  H�  �L  H�      H   ,  �L  FX  �L  G   �  G   �  FX  �L  FX      H   ,  ��  G�  ��  H�  �T  H�  �T  G�  ��  G�      H   ,  �L  E�  �L  FX  �  FX  �  E�  �L  E�      H   ,  �L  J@  �L  K  �  K  �  J@  �L  J@      H   ,  �  G�  �  H�  ��  H�  ��  G�  �  G�      H   ,  ��  G�  ��  H�  ��  H�  ��  G�  ��  G�      H   ,  �L  D�  �L  E�  �  E�  �  D�  �L  D�      H   ,  �L  K�  �L  L�  �  L�  �  K�  �L  K�      H   ,  �L  G�  �L  H�  �  H�  �  G�  �L  G�      H   ,  �L  D   �L  D�  �  D�  �  D   �L  D       H   ,  �,  G�  �,  H�  ��  H�  ��  G�  �,  G�      H   ,  ��  G�  ��  H�  �L  H�  �L  G�  ��  G�      H   ,  �L  Ix  �L  J@  �  J@  �  Ix  �L  Ix      H   ,  ��  G�  ��  H�  ��  H�  ��  G�  ��  G�      H   ,  ��  G�  ��  H�  ��  H�  ��  G�  ��  G�      H   ,  �L  C8  �L  D   �  D   �  C8  �L  C8      H   ,  �L  G   �L  G�  �  G�  �  G   �L  G       H   ,  �L  K  �L  K�  �  K�  �  K  �L  K      H   ,  �L  A�  �L  Bp  �  Bp  �  A�  �L  A�      H   ,  �L  Bp  �L  C8  �  C8  �  Bp  �L  Bp      H   ,  ��  H�  ��  Ix  ��  Ix  ��  H�  ��  H�      H   ,  �  J@  �  K  ��  K  ��  J@  �  J@      H   ,  �  Ix  �  J@  ��  J@  ��  Ix  �  Ix      H   ,  �  H�  �  Ix  ��  Ix  ��  H�  �  H�      H   ,  ��  H�  ��  Ix  �T  Ix  �T  H�  ��  H�      H   ,  ��  K  ��  K�  ��  K�  ��  K  ��  K      H   ,  �,  J@  �,  K  ��  K  ��  J@  �,  J@      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �  K�  �  L�  �d  L�  �d  K�  �  K�      H   ,  ��  K  ��  K�  ��  K�  ��  K  ��  K      H   ,  ��  M`  ��  N(  �L  N(  �L  M`  ��  M`      H   ,  ��  J@  ��  K  ��  K  ��  J@  ��  J@      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  ��  Ix  ��  J@  �L  J@  �L  Ix  ��  Ix      H   ,  �  N(  �  N�  �d  N�  �d  N(  �  N(      H   ,  �,  H�  �,  Ix  ��  Ix  ��  H�  �,  H�      H   ,  �d  L�  �d  M`  �,  M`  �,  L�  �d  L�      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  ��  H�  ��  Ix  ��  Ix  ��  H�  ��  H�      H   ,  ��  J@  ��  K  �L  K  �L  J@  ��  J@      H   ,  �,  N(  �,  N�  ��  N�  ��  N(  �,  N(      H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  �d  J@  �d  K  �,  K  �,  J@  �d  J@      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  ��  K�  ��  L�  �L  L�  �L  K�  ��  K�      H   ,  ~  N(  ~  N�  ~�  N�  ~�  N(  ~  N(      H   ,  �  M`  �  N(  �d  N(  �d  M`  �  M`      H   ,  �,  K�  �,  L�  ��  L�  ��  K�  �,  K�      H   ,  �d  K�  �d  L�  �,  L�  �,  K�  �d  K�      H   ,  ��  H�  ��  Ix  ��  Ix  ��  H�  ��  H�      H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  ��  K  ��  K�  �L  K�  �L  K  ��  K      H   ,  ��  J@  ��  K  ��  K  ��  J@  ��  J@      H   ,  ~�  N(  ~�  N�  �  N�  �  N(  ~�  N(      H   ,  �d  M`  �d  N(  �,  N(  �,  M`  �d  M`      H   ,  �,  M`  �,  N(  ��  N(  ��  M`  �,  M`      H   ,  �,  K  �,  K�  ��  K�  ��  K  �,  K      H   ,  ��  N(  ��  N�  �L  N�  �L  N(  ��  N(      H   ,  �d  Ix  �d  J@  �,  J@  �,  Ix  �d  Ix      H   ,  �d  N(  �d  N�  �,  N�  �,  N(  �d  N(      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �,  L�  �,  M`  ��  M`  ��  L�  �,  L�      H   ,  ~�  M`  ~�  N(  �  N(  �  M`  ~�  M`      H   ,  �  L�  �  M`  �d  M`  �d  L�  �  L�      H   ,  �,  Ix  �,  J@  ��  J@  ��  Ix  �,  Ix      H   ,  ~  M`  ~  N(  ~�  N(  ~�  M`  ~  M`      H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  ��  L�  ��  M`  �L  M`  �L  L�  ��  L�      H   ,  ��  Ix  ��  J@  ��  J@  ��  Ix  ��  Ix      H   ,  ��  H�  ��  Ix  �L  Ix  �L  H�  ��  H�      H   ,  �d  K  �d  K�  �,  K�  �,  K  �d  K      H   ,  ��  Ix  ��  J@  ��  J@  ��  Ix  ��  Ix      H   ,  ��  D�  ��  E�  ��  E�  ��  D�  ��  D�      H   ,  ��  D   ��  D�  �L  D�  �L  D   ��  D       H   ,  ��  E�  ��  FX  ��  FX  ��  E�  ��  E�      H   ,  ��  FX  ��  G   ��  G   ��  FX  ��  FX      H   ,  ��  FX  ��  G   �L  G   �L  FX  ��  FX      H   ,  ��  C8  ��  D   �L  D   �L  C8  ��  C8      H   ,  ��  FX  ��  G   ��  G   ��  FX  ��  FX      H   ,  ��  G   ��  G�  ��  G�  ��  G   ��  G       H   ,  ��  E�  ��  FX  �L  FX  �L  E�  ��  E�      H   ,  ��  G   ��  G�  �L  G�  �L  G   ��  G       H   ,  ��  D�  ��  E�  �L  E�  �L  D�  ��  D�      H   ,  ��  G   ��  G�  ��  G�  ��  G   ��  G       H   ,  ��  G   ��  G�  ��  G�  ��  G   ��  G       H   ,  ��  A�  ��  Bp  ��  Bp  ��  A�  ��  A�      H   ,  ��  FX  ��  G   ��  G   ��  FX  ��  FX      H   ,  �  E�  �  FX  ��  FX  ��  E�  �  E�      H   ,  ��  D   ��  D�  �T  D�  �T  D   ��  D       H   ,  �  D   �  D�  ��  D�  ��  D   �  D       H   ,  ��  D   ��  D�  ��  D�  ��  D   ��  D       H   ,  ��  A�  ��  Bp  �l  Bp  �l  A�  ��  A�      H   ,  ��  E�  ��  FX  ��  FX  ��  E�  ��  E�      H   ,  ��  D   ��  D�  ��  D�  ��  D   ��  D       H   ,  ��  E�  ��  FX  ��  FX  ��  E�  ��  E�      H   ,  �  C8  �  D   ��  D   ��  C8  �  C8      H   ,  �  A�  �  Bp  ��  Bp  ��  A�  �  A�      H   ,  ��  A�  ��  Bp  ��  Bp  ��  A�  ��  A�      H   ,  ��  D�  ��  E�  ��  E�  ��  D�  ��  D�      H   ,  ��  C8  ��  D   �T  D   �T  C8  ��  C8      H   ,  ��  FX  ��  G   �l  G   �l  FX  ��  FX      H   ,  ��  C8  ��  D   ��  D   ��  C8  ��  C8      H   ,  ��  G   ��  G�  �T  G�  �T  G   ��  G       H   ,  �4  Bp  �4  C8  ��  C8  ��  Bp  �4  Bp      H   ,  �l  A�  �l  Bp  �4  Bp  �4  A�  �l  A�      H   ,  ��  D�  ��  E�  �l  E�  �l  D�  ��  D�      H   ,  ��  Bp  ��  C8  �l  C8  �l  Bp  ��  Bp      H   ,  ��  Bp  ��  C8  �T  C8  �T  Bp  ��  Bp      H   ,  ��  C8  ��  D   �l  D   �l  C8  ��  C8      H   ,  ��  C8  ��  D   ��  D   ��  C8  ��  C8      H   ,  �l  D�  �l  E�  �4  E�  �4  D�  �l  D�      H   ,  �  FX  �  G   ��  G   ��  FX  �  FX      H   ,  ��  D�  ��  E�  ��  E�  ��  D�  ��  D�      H   ,  ��  D   ��  D�  ��  D�  ��  D   ��  D       H   ,  ��  C8  ��  D   ��  D   ��  C8  ��  C8      H   ,  ��  E�  ��  FX  �l  FX  �l  E�  ��  E�      H   ,  ��  FX  ��  G   ��  G   ��  FX  ��  FX      H   ,  �4  A�  �4  Bp  ��  Bp  ��  A�  �4  A�      H   ,  ��  A�  ��  Bp  ��  Bp  ��  A�  ��  A�      H   ,  ��  FX  ��  G   �T  G   �T  FX  ��  FX      H   ,  �4  C8  �4  D   ��  D   ��  C8  �4  C8      H   ,  �l  Bp  �l  C8  �4  C8  �4  Bp  �l  Bp      H   ,  �  G   �  G�  ��  G�  ��  G   �  G       H   ,  ��  D�  ��  E�  �T  E�  �T  D�  ��  D�      H   ,  �l  E�  �l  FX  �4  FX  �4  E�  �l  E�      H   ,  �l  C8  �l  D   �4  D   �4  C8  �l  C8      H   ,  ��  Bp  ��  C8  ��  C8  ��  Bp  ��  Bp      H   ,  ��  Bp  ��  C8  ��  C8  ��  Bp  ��  Bp      H   ,  ��  E�  ��  FX  ��  FX  ��  E�  ��  E�      H   ,  ��  D   ��  D�  �l  D�  �l  D   ��  D       H   ,  ��  A�  ��  Bp  �T  Bp  �T  A�  ��  A�      H   ,  �l  D   �l  D�  �4  D�  �4  D   �l  D       H   ,  �  Bp  �  C8  ��  C8  ��  Bp  �  Bp      H   ,  ��  G   ��  G�  �l  G�  �l  G   ��  G       H   ,  ��  Bp  ��  C8  ��  C8  ��  Bp  ��  Bp      H   ,  ��  D�  ��  E�  ��  E�  ��  D�  ��  D�      H   ,  �  D�  �  E�  ��  E�  ��  D�  �  D�      H   ,  ��  E�  ��  FX  �T  FX  �T  E�  ��  E�      H   ,  ��  G   ��  G�  ��  G�  ��  G   ��  G       H   ,  �  K  �  K�  ��  K�  ��  K  �  K      H   ,  �  J@  �  K  ��  K  ��  J@  �  J@      H   ,  �<  N(  �<  N�  �  N�  �  N(  �<  N(      H   ,  �<  G�  �<  H�  �  H�  �  G�  �<  G�      H   ,  �t  K�  �t  L�  �<  L�  �<  K�  �t  K�      H   ,  �<  L�  �<  M`  �  M`  �  L�  �<  L�      H   ,  �  E�  �  FX  ��  FX  ��  E�  �  E�      H   ,  ��  C8  ��  D   ��  D   ��  C8  ��  C8      H   ,  ��  J@  ��  K  ��  K  ��  J@  ��  J@      H   ,  �  J@  �  K  ��  K  ��  J@  �  J@      H   ,  �  G   �  G�  ��  G�  ��  G   �  G       H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �t  G�  �t  H�  �<  H�  �<  G�  �t  G�      H   ,  ��  FX  ��  G   �t  G   �t  FX  ��  FX      H   ,  �  N(  �  N�  ��  N�  ��  N(  �  N(      H   ,  ��  Ix  ��  J@  ��  J@  ��  Ix  ��  Ix      H   ,  �  Ix  �  J@  ��  J@  ��  Ix  �  Ix      H   ,  �<  M`  �<  N(  �  N(  �  M`  �<  M`      H   ,  �t  J@  �t  K  �<  K  �<  J@  �t  J@      H   ,  �  C8  �  D   ��  D   ��  C8  �  C8      H   ,  ��  G   ��  G�  �t  G�  �t  G   ��  G       H   ,  �<  K  �<  K�  �  K�  �  K  �<  K      H   ,  �\  N(  �\  N�  �$  N�  �$  N(  �\  N(      H   ,  ��  H�  ��  Ix  ��  Ix  ��  H�  ��  H�      H   ,  �  Ix  �  J@  ��  J@  ��  Ix  �  Ix      H   ,  ��  K  ��  K�  ��  K�  ��  K  ��  K      H   ,  ��  D   ��  D�  ��  D�  ��  D   ��  D       H   ,  �  FX  �  G   ��  G   ��  FX  �  FX      H   ,  �t  L�  �t  M`  �<  M`  �<  L�  �t  L�      H   ,  ��  E�  ��  FX  �t  FX  �t  E�  ��  E�      H   ,  �t  M`  �t  N(  �<  N(  �<  M`  �t  M`      H   ,  ��  G�  ��  H�  ��  H�  ��  G�  ��  G�      H   ,  ��  M`  ��  N(  ��  N(  ��  M`  ��  M`      H   ,  �  M`  �  N(  ��  N(  ��  M`  �  M`      H   ,  ��  K  ��  K�  �t  K�  �t  K  ��  K      H   ,  �t  G   �t  G�  �<  G�  �<  G   �t  G       H   ,  ��  N(  ��  N�  ��  N�  ��  N(  ��  N(      H   ,  �  K  �  K�  ��  K�  ��  K  �  K      H   ,  �t  FX  �t  G   �<  G   �<  FX  �t  FX      H   ,  ��  G   ��  G�  ��  G�  ��  G   ��  G       H   ,  �  Bp  �  C8  ��  C8  ��  Bp  �  Bp      H   ,  �  H�  �  Ix  ��  Ix  ��  H�  �  H�      H   ,  �t  N(  �t  N�  �<  N�  �<  N(  �t  N(      H   ,  �t  Ix  �t  J@  �<  J@  �<  Ix  �t  Ix      H   ,  �<  J@  �<  K  �  K  �  J@  �<  J@      H   ,  ��  D�  ��  E�  �t  E�  �t  D�  ��  D�      H   ,  �  D   �  D�  ��  D�  ��  D   �  D       H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  ��  FX  ��  G   ��  G   ��  FX  ��  FX      H   ,  �  L�  �  M`  ��  M`  ��  L�  �  L�      H   ,  ��  L�  ��  M`  ��  M`  ��  L�  ��  L�      H   ,  �<  K�  �<  L�  �  L�  �  K�  �<  K�      H   ,  �t  K  �t  K�  �<  K�  �<  K  �t  K      H   ,  ��  Ix  ��  J@  �t  J@  �t  Ix  ��  Ix      H   ,  ��  M`  ��  N(  �t  N(  �t  M`  ��  M`      H   ,  ��  J@  ��  K  �t  K  �t  J@  ��  J@      H   ,  �  D�  �  E�  ��  E�  ��  D�  �  D�      H   ,  ��  E�  ��  FX  ��  FX  ��  E�  ��  E�      H   ,  �<  H�  �<  Ix  �  Ix  �  H�  �<  H�      H   ,  �  K�  �  L�  ��  L�  ��  K�  �  K�      H   ,  �  A�  �  Bp  ��  Bp  ��  A�  �  A�      H   ,  ��  L�  ��  M`  �\  M`  �\  L�  ��  L�      H   ,  ��  K�  ��  L�  ��  L�  ��  K�  ��  K�      H   ,  �t  H�  �t  Ix  �<  Ix  �<  H�  �t  H�      H   ,  �  K�  �  L�  ��  L�  ��  K�  �  K�      H   ,  ��  L�  ��  M`  �t  M`  �t  L�  ��  L�      H   ,  ��  N(  ��  N�  �t  N�  �t  N(  ��  N(      H   ,  ��  D�  ��  E�  ��  E�  ��  D�  ��  D�      H   ,  �  G�  �  H�  ��  H�  ��  G�  �  G�      H   ,  ��  M`  ��  N(  �\  N(  �\  M`  ��  M`      H   ,  ��  N(  ��  N�  �\  N�  �\  N(  ��  N(      H   ,  �<  Ix  �<  J@  �  J@  �  Ix  �<  Ix      H   ,  ��  H�  ��  Ix  �t  Ix  �t  H�  ��  H�      H   ,  ��  K�  ��  L�  �t  L�  �t  K�  ��  K�      H   ,  ��  G�  ��  H�  �t  H�  �t  G�  ��  G�      H   ,  ��  K  ��  K�  ��  K�  ��  K  ��  K      H   ,  �T  @�  �T  A�  �  A�  �  @�  �T  @�      H   ,  �T  @  �T  @�  �  @�  �  @  �T  @      H   ,  �T  ?P  �T  @  �  @  �  ?P  �T  ?P      H   ,  �d  3�  �d  4`  �,  4`  �,  3�  �d  3�      H   ,  �T  =�  �T  >�  �  >�  �  =�  �T  =�      H   ,  �T  <�  �T  =�  �  =�  �  <�  �T  <�      H   ,  �T  <0  �T  <�  �  <�  �  <0  �T  <0      H   ,  �T  ;h  �T  <0  �  <0  �  ;h  �T  ;h      H   ,  �T  :�  �T  ;h  �  ;h  �  :�  �T  :�      H   ,  �T  9�  �T  :�  �  :�  �  9�  �T  9�      H   ,  ��  3�  ��  4`  �L  4`  �L  3�  ��  3�      H   ,  �T  9  �T  9�  �  9�  �  9  �T  9      H   ,  �T  8H  �T  9  �  9  �  8H  �T  8H      H   ,  �T  7�  �T  8H  �  8H  �  7�  �T  7�      H   ,  �T  6�  �T  7�  �  7�  �  6�  �T  6�      H   ,  �  3�  �  4`  ��  4`  ��  3�  �  3�      H   ,  �T  5�  �T  6�  �  6�  �  5�  �T  5�      H   ,  �T  5(  �T  5�  �  5�  �  5(  �T  5(      H   ,  �<  3�  �<  4`  �  4`  �  3�  �<  3�      H   ,  �T  4`  �T  5(  �  5(  �  4`  �T  4`      H   ,  �T  2�  �T  3�  �  3�  �  2�  �T  2�      H   ,  �T  2  �T  2�  �  2�  �  2  �T  2      H   ,  �  3�  �  4`  ��  4`  ��  3�  �  3�      H   ,  �T  1@  �T  2  �  2  �  1@  �T  1@      H   ,  �T  0x  �T  1@  �  1@  �  0x  �T  0x      H   ,  �t  3�  �t  4`  �<  4`  �<  3�  �t  3�      H   ,  �T  /�  �T  0x  �  0x  �  /�  �T  /�      H   ,  �l  3�  �l  4`  �4  4`  �4  3�  �l  3�      H   ,  �L  3�  �L  4`  �  4`  �  3�  �L  3�      H   ,  �T  .�  �T  /�  �  /�  �  .�  �T  .�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  ��  3�  ��  4`  �l  4`  �l  3�  ��  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  ~�  3�  ~�  4`  �  4`  �  3�  ~�  3�      H   ,  �,  3�  �,  4`  ��  4`  ��  3�  �,  3�      H   ,  �  3�  �  4`  �d  4`  �d  3�  �  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  ~  3�  ~  4`  ~�  4`  ~�  3�  ~  3�      H   ,  ��  3�  ��  4`  �t  4`  �t  3�  ��  3�      H   ,  �  3�  �  4`  ��  4`  ��  3�  �  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  �  5(  �  5�  ��  5�  ��  5(  �  5(      H   ,  �  4`  �  5(  ��  5(  ��  4`  �  4`      H   ,  ��  5(  ��  5�  ��  5�  ��  5(  ��  5(      H   ,  �t  5(  �t  5�  �<  5�  �<  5(  �t  5(      H   ,  �  @�  �  A�  ��  A�  ��  @�  �  @�      H   ,  �  :�  �  ;h  ��  ;h  ��  :�  �  :�      H   ,  �t  4`  �t  5(  �<  5(  �<  4`  �t  4`      H   ,  �<  5�  �<  6�  �  6�  �  5�  �<  5�      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  �  <0  �  <�  ��  <�  ��  <0  �  <0      H   ,  �  9�  �  :�  ��  :�  ��  9�  �  9�      H   ,  ��  6�  ��  7�  ��  7�  ��  6�  ��  6�      H   ,  �<  5(  �<  5�  �  5�  �  5(  �<  5(      H   ,  �  9  �  9�  ��  9�  ��  9  �  9      H   ,  �<  4`  �<  5(  �  5(  �  4`  �<  4`      H   ,  ��  9  ��  9�  ��  9�  ��  9  ��  9      H   ,  �t  7�  �t  8H  �<  8H  �<  7�  �t  7�      H   ,  ��  8H  ��  9  ��  9  ��  8H  ��  8H      H   ,  �  8H  �  9  ��  9  ��  8H  �  8H      H   ,  ��  9  ��  9�  �t  9�  �t  9  ��  9      H   ,  ��  5�  ��  6�  ��  6�  ��  5�  ��  5�      H   ,  ��  8H  ��  9  �t  9  �t  8H  ��  8H      H   ,  ��  9�  ��  :�  ��  :�  ��  9�  ��  9�      H   ,  ��  7�  ��  8H  ��  8H  ��  7�  ��  7�      H   ,  ��  7�  ��  8H  �t  8H  �t  7�  ��  7�      H   ,  �  7�  �  8H  ��  8H  ��  7�  �  7�      H   ,  ��  6�  ��  7�  �t  7�  �t  6�  ��  6�      H   ,  ��  5�  ��  6�  �t  6�  �t  5�  ��  5�      H   ,  ��  5(  ��  5�  �t  5�  �t  5(  ��  5(      H   ,  ��  :�  ��  ;h  ��  ;h  ��  :�  ��  :�      H   ,  ��  4`  ��  5(  �t  5(  �t  4`  ��  4`      H   ,  �  ;h  �  <0  ��  <0  ��  ;h  �  ;h      H   ,  �t  6�  �t  7�  �<  7�  �<  6�  �t  6�      H   ,  �  6�  �  7�  ��  7�  ��  6�  �  6�      H   ,  �  5�  �  6�  ��  6�  ��  5�  �  5�      H   ,  �  5(  �  5�  ��  5�  ��  5(  �  5(      H   ,  �  4`  �  5(  ��  5(  ��  4`  �  4`      H   ,  �<  6�  �<  7�  �  7�  �  6�  �<  6�      H   ,  �t  5�  �t  6�  �<  6�  �<  5�  �t  5�      H   ,  �L  9�  �L  :�  �  :�  �  9�  �L  9�      H   ,  �L  9  �L  9�  �  9�  �  9  �L  9      H   ,  �  :�  �  ;h  ��  ;h  ��  :�  �  :�      H   ,  �L  8H  �L  9  �  9  �  8H  �L  8H      H   ,  �4  :�  �4  ;h  ��  ;h  ��  :�  �4  :�      H   ,  �L  7�  �L  8H  �  8H  �  7�  �L  7�      H   ,  �L  6�  �L  7�  �  7�  �  6�  �L  6�      H   ,  �L  5�  �L  6�  �  6�  �  5�  �L  5�      H   ,  �L  5(  �L  5�  �  5�  �  5(  �L  5(      H   ,  �L  4`  �L  5(  �  5(  �  4`  �L  4`      H   ,  ��  :�  ��  ;h  ��  ;h  ��  :�  ��  :�      H   ,  ��  :�  ��  ;h  �l  ;h  �l  :�  ��  :�      H   ,  �l  :�  �l  ;h  �4  ;h  �4  :�  �l  :�      H   ,  ��  :�  ��  ;h  ��  ;h  ��  :�  ��  :�      H   ,  ��  :�  ��  ;h  �T  ;h  �T  :�  ��  :�      H   ,  ��  :�  ��  ;h  ��  ;h  ��  :�  ��  :�      H   ,  �L  :�  �L  ;h  �  ;h  �  :�  �L  :�      H   ,  �l  @�  �l  A�  �4  A�  �4  @�  �l  @�      H   ,  �l  =�  �l  >�  �4  >�  �4  =�  �l  =�      H   ,  ��  <�  ��  =�  ��  =�  ��  <�  ��  <�      H   ,  ��  <0  ��  <�  ��  <�  ��  <0  ��  <0      H   ,  �4  @�  �4  A�  ��  A�  ��  @�  �4  @�      H   ,  �  ;h  �  <0  ��  <0  ��  ;h  �  ;h      H   ,  ��  =�  ��  >�  �T  >�  �T  =�  ��  =�      H   ,  �l  <0  �l  <�  �4  <�  �4  <0  �l  <0      H   ,  ��  >�  ��  ?P  ��  ?P  ��  >�  ��  >�      H   ,  ��  ;h  ��  <0  ��  <0  ��  ;h  ��  ;h      H   ,  �  <0  �  <�  ��  <�  ��  <0  �  <0      H   ,  ��  ;h  ��  <0  �T  <0  �T  ;h  ��  ;h      H   ,  �4  @  �4  @�  ��  @�  ��  @  �4  @      H   ,  ��  @�  ��  A�  �l  A�  �l  @�  ��  @�      H   ,  �4  ;h  �4  <0  ��  <0  ��  ;h  �4  ;h      H   ,  �l  @  �l  @�  �4  @�  �4  @  �l  @      H   ,  ��  >�  ��  ?P  �T  ?P  �T  >�  ��  >�      H   ,  �l  ;h  �l  <0  �4  <0  �4  ;h  �l  ;h      H   ,  ��  @  ��  @�  �l  @�  �l  @  ��  @      H   ,  �4  ?P  �4  @  ��  @  ��  ?P  �4  ?P      H   ,  ��  ?P  ��  @  �l  @  �l  ?P  ��  ?P      H   ,  ��  >�  ��  ?P  �l  ?P  �l  >�  ��  >�      H   ,  �4  >�  �4  ?P  ��  ?P  ��  >�  �4  >�      H   ,  ��  =�  ��  >�  �l  >�  �l  =�  ��  =�      H   ,  ��  @�  ��  A�  ��  A�  ��  @�  ��  @�      H   ,  �l  ?P  �l  @  �4  @  �4  ?P  �l  ?P      H   ,  ��  @  ��  @�  ��  @�  ��  @  ��  @      H   ,  ��  ?P  ��  @  ��  @  ��  ?P  ��  ?P      H   ,  ��  @  ��  @�  ��  @�  ��  @  ��  @      H   ,  ��  >�  ��  ?P  ��  ?P  ��  >�  ��  >�      H   ,  ��  =�  ��  >�  ��  >�  ��  =�  ��  =�      H   ,  ��  <�  ��  =�  �l  =�  �l  <�  ��  <�      H   ,  ��  =�  ��  >�  ��  >�  ��  =�  ��  =�      H   ,  ��  <�  ��  =�  ��  =�  ��  <�  ��  <�      H   ,  ��  <0  ��  <�  ��  <�  ��  <0  ��  <0      H   ,  ��  ;h  ��  <0  ��  <0  ��  ;h  ��  ;h      H   ,  ��  <0  ��  <�  �T  <�  �T  <0  ��  <0      H   ,  �  @�  �  A�  ��  A�  ��  @�  �  @�      H   ,  ��  <0  ��  <�  �l  <�  �l  <0  ��  <0      H   ,  ��  @�  ��  A�  ��  A�  ��  @�  ��  @�      H   ,  ��  @�  ��  A�  �T  A�  �T  @�  ��  @�      H   ,  ��  @  ��  @�  ��  @�  ��  @  ��  @      H   ,  ��  ?P  ��  @  ��  @  ��  ?P  ��  ?P      H   ,  ��  @�  ��  A�  ��  A�  ��  @�  ��  @�      H   ,  ��  >�  ��  ?P  ��  ?P  ��  >�  ��  >�      H   ,  ��  =�  ��  >�  ��  >�  ��  =�  ��  =�      H   ,  �4  =�  �4  >�  ��  >�  ��  =�  �4  =�      H   ,  ��  <�  ��  =�  ��  =�  ��  <�  ��  <�      H   ,  ��  <�  ��  =�  �T  =�  �T  <�  ��  <�      H   ,  ��  @  ��  @�  �T  @�  �T  @  ��  @      H   ,  �4  <0  �4  <�  ��  <�  ��  <0  �4  <0      H   ,  ��  <0  ��  <�  ��  <�  ��  <0  ��  <0      H   ,  ��  ;h  ��  <0  ��  <0  ��  ;h  ��  ;h      H   ,  ��  ;h  ��  <0  �l  <0  �l  ;h  ��  ;h      H   ,  ��  ?P  ��  @  ��  @  ��  ?P  ��  ?P      H   ,  �l  >�  �l  ?P  �4  ?P  �4  >�  �l  >�      H   ,  �l  <�  �l  =�  �4  =�  �4  <�  �l  <�      H   ,  �4  <�  �4  =�  ��  =�  ��  <�  �4  <�      H   ,  ��  ?P  ��  @  �T  @  �T  ?P  ��  ?P      H   ,  �  @  �  @�  ��  @�  ��  @  �  @      H   ,  �  4`  �  5(  �d  5(  �d  4`  �  4`      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  ��  4`  ��  5(  �L  5(  �L  4`  ��  4`      H   ,  ��  5(  ��  5�  ��  5�  ��  5(  ��  5(      H   ,  ~�  4`  ~�  5(  �  5(  �  4`  ~�  4`      H   ,  ��  7�  ��  8H  �L  8H  �L  7�  ��  7�      H   ,  �d  4`  �d  5(  �,  5(  �,  4`  �d  4`      H   ,  ��  5(  ��  5�  �L  5�  �L  5(  ��  5(      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  ��  6�  ��  7�  �L  7�  �L  6�  ��  6�      H   ,  ��  8H  ��  9  �L  9  �L  8H  ��  8H      H   ,  �,  4`  �,  5(  ��  5(  ��  4`  �,  4`      H   ,  ��  5�  ��  6�  �L  6�  �L  5�  ��  5�      H   ,  ~  4`  ~  5(  ~�  5(  ~�  4`  ~  4`      H   ,  ��  5�  ��  6�  ��  6�  ��  5�  ��  5�      H   ,  ��  7�  ��  8H  �T  8H  �T  7�  ��  7�      H   ,  �  5(  �  5�  ��  5�  ��  5(  �  5(      H   ,  �l  9  �l  9�  �4  9�  �4  9  �l  9      H   ,  ��  8H  ��  9  ��  9  ��  8H  ��  8H      H   ,  �4  8H  �4  9  ��  9  ��  8H  �4  8H      H   ,  ��  5(  ��  5�  �l  5�  �l  5(  ��  5(      H   ,  ��  9�  ��  :�  ��  :�  ��  9�  ��  9�      H   ,  �  8H  �  9  ��  9  ��  8H  �  8H      H   ,  ��  6�  ��  7�  �T  7�  �T  6�  ��  6�      H   ,  ��  9  ��  9�  ��  9�  ��  9  ��  9      H   ,  ��  4`  ��  5(  �l  5(  �l  4`  ��  4`      H   ,  ��  5�  ��  6�  �T  6�  �T  5�  ��  5�      H   ,  ��  8H  ��  9  ��  9  ��  8H  ��  8H      H   ,  �  9  �  9�  ��  9�  ��  9  �  9      H   ,  ��  7�  ��  8H  ��  8H  ��  7�  ��  7�      H   ,  ��  9  ��  9�  �T  9�  �T  9  ��  9      H   ,  �  6�  �  7�  ��  7�  ��  6�  �  6�      H   ,  ��  6�  ��  7�  ��  7�  ��  6�  ��  6�      H   ,  ��  6�  ��  7�  �l  7�  �l  6�  ��  6�      H   ,  ��  5�  ��  6�  ��  6�  ��  5�  ��  5�      H   ,  ��  9�  ��  :�  ��  :�  ��  9�  ��  9�      H   ,  �l  5�  �l  6�  �4  6�  �4  5�  �l  5�      H   ,  �l  8H  �l  9  �4  9  �4  8H  �l  8H      H   ,  �l  7�  �l  8H  �4  8H  �4  7�  �l  7�      H   ,  ��  5(  ��  5�  ��  5�  ��  5(  ��  5(      H   ,  ��  7�  ��  8H  �l  8H  �l  7�  ��  7�      H   ,  ��  9�  ��  :�  �T  :�  �T  9�  ��  9�      H   ,  �4  9  �4  9�  ��  9�  ��  9  �4  9      H   ,  �  5�  �  6�  ��  6�  ��  5�  �  5�      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  ��  8H  ��  9  �T  9  �T  8H  ��  8H      H   ,  �l  9�  �l  :�  �4  :�  �4  9�  �l  9�      H   ,  ��  9  ��  9�  ��  9�  ��  9  ��  9      H   ,  �  9�  �  :�  ��  :�  ��  9�  �  9�      H   ,  �  4`  �  5(  ��  5(  ��  4`  �  4`      H   ,  ��  9�  ��  :�  �l  :�  �l  9�  ��  9�      H   ,  ��  9�  ��  :�  ��  :�  ��  9�  ��  9�      H   ,  �  7�  �  8H  ��  8H  ��  7�  �  7�      H   ,  ��  9  ��  9�  ��  9�  ��  9  ��  9      H   ,  ��  9  ��  9�  �l  9�  �l  9  ��  9      H   ,  ��  8H  ��  9  ��  9  ��  8H  ��  8H      H   ,  ��  5�  ��  6�  �l  6�  �l  5�  ��  5�      H   ,  ��  7�  ��  8H  ��  8H  ��  7�  ��  7�      H   ,  �4  9�  �4  :�  ��  :�  ��  9�  �4  9�      H   ,  ��  8H  ��  9  �l  9  �l  8H  ��  8H      H   ,  �l  6�  �l  7�  �4  7�  �4  6�  �l  6�      H   ,  ��  6�  ��  7�  ��  7�  ��  6�  ��  6�      H   ,  �L  0x  �L  1@  �  1@  �  0x  �L  0x      H   ,  �L  /�  �L  0x  �  0x  �  /�  �L  /�      H   ,  �L  .�  �L  /�  �  /�  �  .�  �L  .�      H   ,  �L  .   �L  .�  �  .�  �  .   �L  .       H   ,  �L  -X  �L  .   �  .   �  -X  �L  -X      H   ,  �L  ,�  �L  -X  �  -X  �  ,�  �L  ,�      H   ,  ��  ,�  ��  -X  ��  -X  ��  ,�  ��  ,�      H   ,  �d  ,�  �d  -X  �,  -X  �,  ,�  �d  ,�      H   ,  ��  ,�  ��  -X  ��  -X  ��  ,�  ��  ,�      H   ,  ��  ,�  ��  -X  �L  -X  �L  ,�  ��  ,�      H   ,  �L  2�  �L  3�  �  3�  �  2�  �L  2�      H   ,  �,  ,�  �,  -X  ��  -X  ��  ,�  �,  ,�      H   ,  �L  2  �L  2�  �  2�  �  2  �L  2      H   ,  �  ,�  �  -X  �d  -X  �d  ,�  �  ,�      H   ,  �L  1@  �L  2  �  2  �  1@  �L  1@      H   ,  ��  1@  ��  2  �T  2  �T  1@  ��  1@      H   ,  ��  2  ��  2�  �l  2�  �l  2  ��  2      H   ,  ��  0x  ��  1@  �T  1@  �T  0x  ��  0x      H   ,  ��  1@  ��  2  �l  2  �l  1@  ��  1@      H   ,  ��  /�  ��  0x  �T  0x  �T  /�  ��  /�      H   ,  �  2  �  2�  ��  2�  ��  2  �  2      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  .�  ��  /�  �T  /�  �T  .�  ��  .�      H   ,  ��  0x  ��  1@  �l  1@  �l  0x  ��  0x      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  �  1@  �  2  ��  2  ��  1@  �  1@      H   ,  ��  /�  ��  0x  �l  0x  �l  /�  ��  /�      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  �4  2�  �4  3�  ��  3�  ��  2�  �4  2�      H   ,  �l  .�  �l  /�  �4  /�  �4  .�  �l  .�      H   ,  �l  /�  �l  0x  �4  0x  �4  /�  �l  /�      H   ,  �  0x  �  1@  ��  1@  ��  0x  �  0x      H   ,  ��  .�  ��  /�  �l  /�  �l  .�  ��  .�      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �4  2  �4  2�  ��  2�  ��  2  �4  2      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �4  1@  �4  2  ��  2  ��  1@  �4  1@      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �l  2�  �l  3�  �4  3�  �4  2�  �l  2�      H   ,  �  /�  �  0x  ��  0x  ��  /�  �  /�      H   ,  ��  2  ��  2�  �T  2�  �T  2  ��  2      H   ,  �4  0x  �4  1@  ��  1@  ��  0x  �4  0x      H   ,  �  2�  �  3�  ��  3�  ��  2�  �  2�      H   ,  �l  2  �l  2�  �4  2�  �4  2  �l  2      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  �  .�  �  /�  ��  /�  ��  .�  �  .�      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  �l  0x  �l  1@  �4  1@  �4  0x  �l  0x      H   ,  �4  /�  �4  0x  ��  0x  ��  /�  �4  /�      H   ,  ��  2�  ��  3�  �l  3�  �l  2�  ��  2�      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �l  1@  �l  2  �4  2  �4  1@  �l  1@      H   ,  ��  2�  ��  3�  �T  3�  �T  2�  ��  2�      H   ,  �4  .�  �4  /�  ��  /�  ��  .�  �4  .�      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  �d  1@  �d  2  �,  2  �,  1@  �d  1@      H   ,  �,  0x  �,  1@  ��  1@  ��  0x  �,  0x      H   ,  ��  0x  ��  1@  �L  1@  �L  0x  ��  0x      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  �d  2  �d  2�  �,  2�  �,  2  �d  2      H   ,  ��  -X  ��  .   �L  .   �L  -X  ��  -X      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  �,  /�  �,  0x  ��  0x  ��  /�  �,  /�      H   ,  ��  .�  ��  /�  �L  /�  �L  .�  ��  .�      H   ,  �d  .�  �d  /�  �,  /�  �,  .�  �d  .�      H   ,  �,  .�  �,  /�  ��  /�  ��  .�  �,  .�      H   ,  ~  0x  ~  1@  ~�  1@  ~�  0x  ~  0x      H   ,  ~  1@  ~  2  ~�  2  ~�  1@  ~  1@      H   ,  �,  .   �,  .�  ��  .�  ��  .   �,  .       H   ,  �d  2�  �d  3�  �,  3�  �,  2�  �d  2�      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �d  .   �d  .�  �,  .�  �,  .   �d  .       H   ,  �,  -X  �,  .   ��  .   ��  -X  �,  -X      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  2  ��  2�  �L  2�  �L  2  ��  2      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  ��  -X  ��  .   ��  .   ��  -X  ��  -X      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ~�  2�  ~�  3�  �  3�  �  2�  ~�  2�      H   ,  �  2�  �  3�  �d  3�  �d  2�  �  2�      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �  2  �  2�  �d  2�  �d  2  �  2      H   ,  ��  1@  ��  2  �L  2  �L  1@  ��  1@      H   ,  �  1@  �  2  �d  2  �d  1@  �  1@      H   ,  ~�  2  ~�  2�  �  2�  �  2  ~�  2      H   ,  ��  2�  ��  3�  �L  3�  �L  2�  ��  2�      H   ,  ��  -X  ��  .   ��  .   ��  -X  ��  -X      H   ,  �  0x  �  1@  �d  1@  �d  0x  �  0x      H   ,  ��  .   ��  .�  �L  .�  �L  .   ��  .       H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ~�  1@  ~�  2  �  2  �  1@  ~�  1@      H   ,  �,  2�  �,  3�  ��  3�  ��  2�  �,  2�      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �d  -X  �d  .   �,  .   �,  -X  �d  -X      H   ,  ��  /�  ��  0x  �L  0x  �L  /�  ��  /�      H   ,  ~  2�  ~  3�  ~�  3�  ~�  2�  ~  2�      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ~�  0x  ~�  1@  �  1@  �  0x  ~�  0x      H   ,  �,  2  �,  2�  ��  2�  ��  2  �,  2      H   ,  �d  /�  �d  0x  �,  0x  �,  /�  �d  /�      H   ,  �,  1@  �,  2  ��  2  ��  1@  �,  1@      H   ,  �d  0x  �d  1@  �,  1@  �,  0x  �d  0x      H   ,  ~  2  ~  2�  ~�  2�  ~�  2  ~  2      H   ,  �d  (�  �d  )p  �,  )p  �,  (�  �d  (�      H   ,  ��  &P  ��  '  ��  '  ��  &P  ��  &P      H   ,  ~  '  ~  '�  ~�  '�  ~�  '  ~  '      H   ,  ��  *8  ��  +   ��  +   ��  *8  ��  *8      H   ,  �d  &P  �d  '  �,  '  �,  &P  �d  &P      H   ,  �  '�  �  (�  �d  (�  �d  '�  �  '�      H   ,  �d  +   �d  +�  �,  +�  �,  +   �d  +       H   ,  ��  *8  ��  +   �L  +   �L  *8  ��  *8      H   ,  �d  '�  �d  (�  �,  (�  �,  '�  �d  '�      H   ,  �d  )p  �d  *8  �,  *8  �,  )p  �d  )p      H   ,  ~�  (�  ~�  )p  �  )p  �  (�  ~�  (�      H   ,  ��  +�  ��  ,�  �L  ,�  �L  +�  ��  +�      H   ,  ��  )p  ��  *8  ��  *8  ��  )p  ��  )p      H   ,  ��  '�  ��  (�  ��  (�  ��  '�  ��  '�      H   ,  �,  '  �,  '�  ��  '�  ��  '  �,  '      H   ,  �  (�  �  )p  �d  )p  �d  (�  �  (�      H   ,  �,  +�  �,  ,�  ��  ,�  ��  +�  �,  +�      H   ,  ��  +   ��  +�  ��  +�  ��  +   ��  +       H   ,  �,  &P  �,  '  ��  '  ��  &P  �,  &P      H   ,  ��  )p  ��  *8  ��  *8  ��  )p  ��  )p      H   ,  ��  (�  ��  )p  ��  )p  ��  (�  ��  (�      H   ,  ��  +�  ��  ,�  ��  ,�  ��  +�  ��  +�      H   ,  �d  +�  �d  ,�  �,  ,�  �,  +�  �d  +�      H   ,  ~�  '�  ~�  (�  �  (�  �  '�  ~�  '�      H   ,  �  '  �  '�  �d  '�  �d  '  �  '      H   ,  ~�  *8  ~�  +   �  +   �  *8  ~�  *8      H   ,  ��  '�  ��  (�  ��  (�  ��  '�  ��  '�      H   ,  �,  +   �,  +�  ��  +�  ��  +   �,  +       H   ,  ��  (�  ��  )p  ��  )p  ��  (�  ��  (�      H   ,  ��  *8  ��  +   ��  +   ��  *8  ��  *8      H   ,  ~�  '  ~�  '�  �  '�  �  '  ~�  '      H   ,  ��  +   ��  +�  ��  +�  ��  +   ��  +       H   ,  �d  '  �d  '�  �,  '�  �,  '  �d  '      H   ,  �  +�  �  ,�  �d  ,�  �d  +�  �  +�      H   ,  �d  *8  �d  +   �,  +   �,  *8  �d  *8      H   ,  ��  +   ��  +�  �L  +�  �L  +   ��  +       H   ,  ��  '  ��  '�  ��  '�  ��  '  ��  '      H   ,  �,  '�  �,  (�  ��  (�  ��  '�  �,  '�      H   ,  �,  *8  �,  +   ��  +   ��  *8  �,  *8      H   ,  �,  (�  �,  )p  ��  )p  ��  (�  �,  (�      H   ,  ~  &P  ~  '  ~�  '  ~�  &P  ~  &P      H   ,  �  +   �  +�  �d  +�  �d  +   �  +       H   ,  ~�  )p  ~�  *8  �  *8  �  )p  ~�  )p      H   ,  �  &P  �  '  �d  '  �d  &P  �  &P      H   ,  �  *8  �  +   �d  +   �d  *8  �  *8      H   ,  ~�  &P  ~�  '  �  '  �  &P  ~�  &P      H   ,  �,  )p  �,  *8  ��  *8  ��  )p  �,  )p      H   ,  �  )p  �  *8  �d  *8  �d  )p  �  )p      H   ,  ��  '  ��  '�  ��  '�  ��  '  ��  '      H   ,  ��  +�  ��  ,�  ��  ,�  ��  +�  ��  +�      H   ,  �\  (�  �\  )p  �$  )p  �$  (�  �\  (�      H   ,  �\  )p  �\  *8  �$  *8  �$  )p  �\  )p      H   ,  ��  ,�  ��  -X  �|  -X  �|  ,�  ��  ,�      H   ,  �\  2  �\  2�  �$  2�  �$  2  �\  2      H   ,  �\  1@  �\  2  �$  2  �$  1@  �\  1@      H   ,  �\  0x  �\  1@  �$  1@  �$  0x  �\  0x      H   ,  �\  /�  �\  0x  �$  0x  �$  /�  �\  /�      H   ,  �\  *8  �\  +   �$  +   �$  *8  �\  *8      H   ,  �\  .�  �\  /�  �$  /�  �$  .�  �\  .�      H   ,  �\  .   �\  .�  �$  .�  �$  .   �\  .       H   ,  �\  -X  �\  .   �$  .   �$  -X  �\  -X      H   ,  �\  ,�  �\  -X  �$  -X  �$  ,�  �\  ,�      H   ,  �|  ,�  �|  -X  �D  -X  �D  ,�  �|  ,�      H   ,  �  ,�  �  -X  ��  -X  ��  ,�  �  ,�      H   ,  �$  ,�  �$  -X  ��  -X  ��  ,�  �$  ,�      H   ,  �\  +�  �\  ,�  �$  ,�  �$  +�  �\  +�      H   ,  ��  ,�  ��  -X  ��  -X  ��  ,�  ��  ,�      H   ,  ��  ,�  ��  -X  �\  -X  �\  ,�  ��  ,�      H   ,  ��  ,�  ��  -X  ��  -X  ��  ,�  ��  ,�      H   ,  �\  +   �\  +�  �$  +�  �$  +   �\  +       H   ,  ��  /�  ��  0x  �d  0x  �d  /�  ��  /�      H   ,  �  /�  �  0x  ��  0x  ��  /�  �  /�      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  �D  .�  �D  /�  �  /�  �  .�  �D  .�      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  �D  .   �D  .�  �  .�  �  .   �D  .       H   ,  ��  2  ��  2�  �d  2�  �d  2  ��  2      H   ,  ��  .�  ��  /�  �d  /�  �d  .�  ��  .�      H   ,  �D  2  �D  2�  �  2�  �  2  �D  2      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  �  1@  �  2  ��  2  ��  1@  �  1@      H   ,  ��  2  ��  2�  �|  2�  �|  2  ��  2      H   ,  ��  .   ��  .�  �d  .�  �d  .   ��  .       H   ,  �  .   �  .�  ��  .�  ��  .   �  .       H   ,  ��  .�  ��  /�  �|  /�  �|  .�  ��  .�      H   ,  �|  2  �|  2�  �D  2�  �D  2  �|  2      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  .   ��  .�  �|  .�  �|  .   ��  .       H   ,  �|  1@  �|  2  �D  2  �D  1@  �|  1@      H   ,  �$  2  �$  2�  ��  2�  ��  2  �$  2      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  �|  0x  �|  1@  �D  1@  �D  0x  �|  0x      H   ,  ��  -X  ��  .   �|  .   �|  -X  ��  -X      H   ,  ��  0x  ��  1@  �|  1@  �|  0x  ��  0x      H   ,  �$  1@  �$  2  ��  2  ��  1@  �$  1@      H   ,  �|  /�  �|  0x  �D  0x  �D  /�  �|  /�      H   ,  �$  0x  �$  1@  ��  1@  ��  0x  �$  0x      H   ,  ��  -X  ��  .   ��  .   ��  -X  ��  -X      H   ,  ��  1@  ��  2  �d  2  �d  1@  ��  1@      H   ,  �$  /�  �$  0x  ��  0x  ��  /�  �$  /�      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �|  .�  �|  /�  �D  /�  �D  .�  �|  .�      H   ,  �$  .�  �$  /�  ��  /�  ��  .�  �$  .�      H   ,  �|  .   �|  .�  �D  .�  �D  .   �|  .       H   ,  �$  .   �$  .�  ��  .�  ��  .   �$  .       H   ,  �  0x  �  1@  ��  1@  ��  0x  �  0x      H   ,  ��  /�  ��  0x  �|  0x  �|  /�  ��  /�      H   ,  �$  -X  �$  .   ��  .   ��  -X  �$  -X      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �D  1@  �D  2  �  2  �  1@  �D  1@      H   ,  �  2  �  2�  ��  2�  ��  2  �  2      H   ,  ��  0x  ��  1@  �d  1@  �d  0x  ��  0x      H   ,  �  .�  �  /�  ��  /�  ��  .�  �  .�      H   ,  ��  1@  ��  2  �|  2  �|  1@  ��  1@      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �D  0x  �D  1@  �  1@  �  0x  �D  0x      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �D  /�  �D  0x  �  0x  �  /�  �D  /�      H   ,  �<  2�  �<  3�  �  3�  �  2�  �<  2�      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  �t  1@  �t  2  �<  2  �<  1@  �t  1@      H   ,  �t  2  �t  2�  �<  2�  �<  2  �t  2      H   ,  ��  .�  ��  /�  �t  /�  �t  .�  ��  .�      H   ,  ��  /�  ��  0x  �t  0x  �t  /�  ��  /�      H   ,  �  1@  �  2  ��  2  ��  1@  �  1@      H   ,  �t  /�  �t  0x  �<  0x  �<  /�  �t  /�      H   ,  ��  .�  ��  /�  �\  /�  �\  .�  ��  .�      H   ,  �  0x  �  1@  ��  1@  ��  0x  �  0x      H   ,  �  -X  �  .   ��  .   ��  -X  �  -X      H   ,  ��  1@  ��  2  �\  2  �\  1@  ��  1@      H   ,  �  .�  �  /�  ��  /�  ��  .�  �  .�      H   ,  �  2�  �  3�  ��  3�  ��  2�  �  2�      H   ,  �<  .   �<  .�  �  .�  �  .   �<  .       H   ,  �<  /�  �<  0x  �  0x  �  /�  �<  /�      H   ,  ��  .   ��  .�  �t  .�  �t  .   ��  .       H   ,  ��  2�  ��  3�  �\  3�  �\  2�  ��  2�      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �<  1@  �<  2  �  2  �  1@  �<  1@      H   ,  ��  -X  ��  .   ��  .   ��  -X  ��  -X      H   ,  ��  .   ��  .�  �\  .�  �\  .   ��  .       H   ,  �t  .�  �t  /�  �<  /�  �<  .�  �t  .�      H   ,  �<  0x  �<  1@  �  1@  �  0x  �<  0x      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  0x  ��  1@  �\  1@  �\  0x  ��  0x      H   ,  ��  2  ��  2�  �t  2�  �t  2  ��  2      H   ,  �<  2  �<  2�  �  2�  �  2  �<  2      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �  0x  �  1@  ��  1@  ��  0x  �  0x      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  0x  ��  1@  �t  1@  �t  0x  ��  0x      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  -X  ��  .   �\  .   �\  -X  ��  -X      H   ,  �  2  �  2�  ��  2�  ��  2  �  2      H   ,  �t  .   �t  .�  �<  .�  �<  .   �t  .       H   ,  �<  -X  �<  .   �  .   �  -X  �<  -X      H   ,  �  .�  �  /�  ��  /�  ��  .�  �  .�      H   ,  �t  2�  �t  3�  �<  3�  �<  2�  �t  2�      H   ,  �t  0x  �t  1@  �<  1@  �<  0x  �t  0x      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  �<  .�  �<  /�  �  /�  �  .�  �<  .�      H   ,  ��  2  ��  2�  �\  2�  �\  2  ��  2      H   ,  �  2�  �  3�  ��  3�  ��  2�  �  2�      H   ,  ��  2�  ��  3�  �t  3�  �t  2�  ��  2�      H   ,  �  .   �  .�  ��  .�  ��  .   �  .       H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �  2  �  2�  ��  2�  ��  2  �  2      H   ,  ��  /�  ��  0x  �\  0x  �\  /�  ��  /�      H   ,  �  /�  �  0x  ��  0x  ��  /�  �  /�      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  ��  1@  ��  2  �t  2  �t  1@  ��  1@      H   ,  �  1@  �  2  ��  2  ��  1@  �  1@      H   ,  �  /�  �  0x  ��  0x  ��  /�  �  /�      H   ,  ��  +   ��  +�  �\  +�  �\  +   ��  +       H   ,  ��  +�  ��  ,�  ��  ,�  ��  +�  ��  +�      H   ,  ��  *8  ��  +   �\  +   �\  *8  ��  *8      H   ,  ��  +�  ��  ,�  �\  ,�  �\  +�  ��  +�      H   ,  ��  +   ��  +�  ��  +�  ��  +   ��  +       H   ,  �D  +   �D  +�  �  +�  �  +   �D  +       H   ,  ��  (�  ��  )p  �|  )p  �|  (�  ��  (�      H   ,  ��  +�  ��  ,�  �|  ,�  �|  +�  ��  +�      H   ,  �$  *8  �$  +   ��  +   ��  *8  �$  *8      H   ,  ��  '�  ��  (�  ��  (�  ��  '�  ��  '�      H   ,  �|  &P  �|  '  �D  '  �D  &P  �|  &P      H   ,  �  '�  �  (�  ��  (�  ��  '�  �  '�      H   ,  ��  '  ��  '�  �d  '�  �d  '  ��  '      H   ,  �|  '�  �|  (�  �D  (�  �D  '�  �|  '�      H   ,  ��  )p  ��  *8  ��  *8  ��  )p  ��  )p      H   ,  �$  )p  �$  *8  ��  *8  ��  )p  �$  )p      H   ,  �  (�  �  )p  ��  )p  ��  (�  �  (�      H   ,  ��  *8  ��  +   ��  +   ��  *8  ��  *8      H   ,  �  )p  �  *8  ��  *8  ��  )p  �  )p      H   ,  ��  (�  ��  )p  ��  )p  ��  (�  ��  (�      H   ,  �|  )p  �|  *8  �D  *8  �D  )p  �|  )p      H   ,  �D  *8  �D  +   �  +   �  *8  �D  *8      H   ,  �  &P  �  '  ��  '  ��  &P  �  &P      H   ,  �|  (�  �|  )p  �D  )p  �D  (�  �|  (�      H   ,  ��  &P  ��  '  ��  '  ��  &P  ��  &P      H   ,  �$  '�  �$  (�  ��  (�  ��  '�  �$  '�      H   ,  ��  )p  ��  *8  �|  *8  �|  )p  ��  )p      H   ,  �D  )p  �D  *8  �  *8  �  )p  �D  )p      H   ,  ��  '  ��  '�  ��  '�  ��  '  ��  '      H   ,  ��  &P  ��  '  �d  '  �d  &P  ��  &P      H   ,  �D  (�  �D  )p  �  )p  �  (�  �D  (�      H   ,  ��  '  ��  '�  �|  '�  �|  '  ��  '      H   ,  �$  +   �$  +�  ��  +�  ��  +   �$  +       H   ,  �D  '�  �D  (�  �  (�  �  '�  �D  '�      H   ,  ��  '�  ��  (�  ��  (�  ��  '�  ��  '�      H   ,  �|  '  �|  '�  �D  '�  �D  '  �|  '      H   ,  �|  +�  �|  ,�  �D  ,�  �D  +�  �|  +�      H   ,  ��  +�  ��  ,�  ��  ,�  ��  +�  ��  +�      H   ,  �D  '  �D  '�  �  '�  �  '  �D  '      H   ,  �|  *8  �|  +   �D  +   �D  *8  �|  *8      H   ,  ��  *8  ��  +   �|  +   �|  *8  ��  *8      H   ,  �$  +�  �$  ,�  ��  ,�  ��  +�  �$  +�      H   ,  ��  +   ��  +�  ��  +�  ��  +   ��  +       H   ,  ��  +   ��  +�  �|  +�  �|  +   ��  +       H   ,  �|  +   �|  +�  �D  +�  �D  +   �|  +       H   ,  ��  '  ��  '�  ��  '�  ��  '  ��  '      H   ,  ��  &P  ��  '  ��  '  ��  &P  ��  &P      H   ,  ��  '�  ��  (�  �d  (�  �d  '�  ��  '�      H   ,  �$  (�  �$  )p  ��  )p  ��  (�  �$  (�      H   ,  �D  &P  �D  '  �  '  �  &P  �D  &P      H   ,  ��  '�  ��  (�  �|  (�  �|  '�  ��  '�      H   ,  ��  (�  ��  )p  ��  )p  ��  (�  ��  (�      H   ,  �  *8  �  +   ��  +   ��  *8  �  *8      H   ,  �  '  �  '�  ��  '�  ��  '  �  '      H   ,  ��  &P  ��  '  �|  '  �|  &P  ��  &P      H   ,  x�  3�  x�  4`  y\  4`  y\  3�  x�  3�      H   ,  s  3�  s  4`  s�  4`  s�  3�  s  3�      H   ,  o�  9  o�  9�  p�  9�  p�  9  o�  9      H   ,  v<  3�  v<  4`  w  4`  w  3�  v<  3�      H   ,  rT  3�  rT  4`  s  4`  s  3�  rT  3�      H   ,  o�  8H  o�  9  p�  9  p�  8H  o�  8H      H   ,  z�  3�  z�  4`  {�  4`  {�  3�  z�  3�      H   ,  p�  3�  p�  4`  q�  4`  q�  3�  p�  3�      H   ,  ut  3�  ut  4`  v<  4`  v<  3�  ut  3�      H   ,  o�  7�  o�  8H  p�  8H  p�  7�  o�  7�      H   ,  z$  3�  z$  4`  z�  4`  z�  3�  z$  3�      H   ,  o�  6�  o�  7�  p�  7�  p�  6�  o�  6�      H   ,  o�  5�  o�  6�  p�  6�  p�  5�  o�  5�      H   ,  w�  3�  w�  4`  x�  4`  x�  3�  w�  3�      H   ,  o�  5(  o�  5�  p�  5�  p�  5(  o�  5(      H   ,  o�  4`  o�  5(  p�  5(  p�  4`  o�  4`      H   ,  q�  3�  q�  4`  rT  4`  rT  3�  q�  3�      H   ,  s�  3�  s�  4`  t�  4`  t�  3�  s�  3�      H   ,  w  3�  w  4`  w�  4`  w�  3�  w  3�      H   ,  y\  3�  y\  4`  z$  4`  z$  3�  y\  3�      H   ,  t�  3�  t�  4`  ut  4`  ut  3�  t�  3�      H   ,  {�  3�  {�  4`  ||  4`  ||  3�  {�  3�      H   ,  ||  3�  ||  4`  }D  4`  }D  3�  ||  3�      H   ,  }D  3�  }D  4`  ~  4`  ~  3�  }D  3�      H   ,  z�  5(  z�  5�  {�  5�  {�  5(  z�  5(      H   ,  p�  5�  p�  6�  q�  6�  q�  5�  p�  5�      H   ,  ut  5(  ut  5�  v<  5�  v<  5(  ut  5(      H   ,  rT  6�  rT  7�  s  7�  s  6�  rT  6�      H   ,  v<  4`  v<  5(  w  5(  w  4`  v<  4`      H   ,  z�  4`  z�  5(  {�  5(  {�  4`  z�  4`      H   ,  {�  4`  {�  5(  ||  5(  ||  4`  {�  4`      H   ,  {�  5(  {�  5�  ||  5�  ||  5(  {�  5(      H   ,  s  7�  s  8H  s�  8H  s�  7�  s  7�      H   ,  ut  6�  ut  7�  v<  7�  v<  6�  ut  6�      H   ,  z$  5(  z$  5�  z�  5�  z�  5(  z$  5(      H   ,  p�  5(  p�  5�  q�  5�  q�  5(  p�  5(      H   ,  x�  4`  x�  5(  y\  5(  y\  4`  x�  4`      H   ,  s�  7�  s�  8H  t�  8H  t�  7�  s�  7�      H   ,  ||  4`  ||  5(  }D  5(  }D  4`  ||  4`      H   ,  x�  5(  x�  5�  y\  5�  y\  5(  x�  5(      H   ,  v<  5(  v<  5�  w  5�  w  5(  v<  5(      H   ,  s�  6�  s�  7�  t�  7�  t�  6�  s�  6�      H   ,  s�  5�  s�  6�  t�  6�  t�  5�  s�  5�      H   ,  p�  6�  p�  7�  q�  7�  q�  6�  p�  6�      H   ,  w  5�  w  6�  w�  6�  w�  5�  w  5�      H   ,  s�  5(  s�  5�  t�  5�  t�  5(  s�  5(      H   ,  s  6�  s  7�  s�  7�  s�  6�  s  6�      H   ,  s�  4`  s�  5(  t�  5(  t�  4`  s�  4`      H   ,  x�  5�  x�  6�  y\  6�  y\  5�  x�  5�      H   ,  q�  8H  q�  9  rT  9  rT  8H  q�  8H      H   ,  rT  4`  rT  5(  s  5(  s  4`  rT  4`      H   ,  y\  5�  y\  6�  z$  6�  z$  5�  y\  5�      H   ,  rT  5�  rT  6�  s  6�  s  5�  rT  5�      H   ,  t�  6�  t�  7�  ut  7�  ut  6�  t�  6�      H   ,  w  4`  w  5(  w�  5(  w�  4`  w  4`      H   ,  y\  5(  y\  5�  z$  5�  z$  5(  y\  5(      H   ,  q�  7�  q�  8H  rT  8H  rT  7�  q�  7�      H   ,  t�  5�  t�  6�  ut  6�  ut  5�  t�  5�      H   ,  ut  4`  ut  5(  v<  5(  v<  4`  ut  4`      H   ,  y\  4`  y\  5(  z$  5(  z$  4`  y\  4`      H   ,  t�  5(  t�  5�  ut  5�  ut  5(  t�  5(      H   ,  s  5�  s  6�  s�  6�  s�  5�  s  5�      H   ,  q�  6�  q�  7�  rT  7�  rT  6�  q�  6�      H   ,  t�  4`  t�  5(  ut  5(  ut  4`  t�  4`      H   ,  w  6�  w  7�  w�  7�  w�  6�  w  6�      H   ,  w�  5�  w�  6�  x�  6�  x�  5�  w�  5�      H   ,  v<  6�  v<  7�  w  7�  w  6�  v<  6�      H   ,  p�  4`  p�  5(  q�  5(  q�  4`  p�  4`      H   ,  rT  5(  rT  5�  s  5�  s  5(  rT  5(      H   ,  w�  5(  w�  5�  x�  5�  x�  5(  w�  5(      H   ,  q�  5�  q�  6�  rT  6�  rT  5�  q�  5�      H   ,  }D  5(  }D  5�  ~  5�  ~  5(  }D  5(      H   ,  s  5(  s  5�  s�  5�  s�  5(  s  5(      H   ,  ut  5�  ut  6�  v<  6�  v<  5�  ut  5�      H   ,  rT  7�  rT  8H  s  8H  s  7�  rT  7�      H   ,  z$  4`  z$  5(  z�  5(  z�  4`  z$  4`      H   ,  }D  4`  }D  5(  ~  5(  ~  4`  }D  4`      H   ,  w  5(  w  5�  w�  5�  w�  5(  w  5(      H   ,  q�  5(  q�  5�  rT  5�  rT  5(  q�  5(      H   ,  w�  4`  w�  5(  x�  5(  x�  4`  w�  4`      H   ,  p�  8H  p�  9  q�  9  q�  8H  p�  8H      H   ,  ||  5(  ||  5�  }D  5�  }D  5(  ||  5(      H   ,  p�  7�  p�  8H  q�  8H  q�  7�  p�  7�      H   ,  s  4`  s  5(  s�  5(  s�  4`  s  4`      H   ,  q�  4`  q�  5(  rT  5(  rT  4`  q�  4`      H   ,  v<  5�  v<  6�  w  6�  w  5�  v<  5�      H   ,  h�  7�  h�  8H  i�  8H  i�  7�  h�  7�      H   ,  h�  9  h�  9�  i�  9�  i�  9  h�  9      H   ,  h�  9�  h�  :�  i�  :�  i�  9�  h�  9�      H   ,  j�  :�  j�  ;h  kL  ;h  kL  :�  j�  :�      H   ,  i�  :�  i�  ;h  j�  ;h  j�  :�  i�  :�      H   ,  h,  :�  h,  ;h  h�  ;h  h�  :�  h,  :�      H   ,  f�  :�  f�  ;h  gd  ;h  gd  :�  f�  :�      H   ,  e  :�  e  ;h  e�  ;h  e�  :�  e  :�      H   ,  h�  8H  h�  9  i�  9  i�  8H  h�  8H      H   ,  h�  ;h  h�  <0  i�  <0  i�  ;h  h�  ;h      H   ,  h�  :�  h�  ;h  i�  ;h  i�  :�  h�  :�      H   ,  l  :�  l  ;h  l�  ;h  l�  :�  l  :�      H   ,  gd  :�  gd  ;h  h,  ;h  h,  :�  gd  :�      H   ,  h�  <0  h�  <�  i�  <�  i�  <0  h�  <0      H   ,  kL  :�  kL  ;h  l  ;h  l  :�  kL  :�      H   ,  e�  :�  e�  ;h  f�  ;h  f�  :�  e�  :�      H   ,  h�  <�  h�  =�  i�  =�  i�  <�  h�  <�      H   ,  i�  <0  i�  <�  j�  <�  j�  <0  i�  <0      H   ,  kL  ;h  kL  <0  l  <0  l  ;h  kL  ;h      H   ,  i�  ;h  i�  <0  j�  <0  j�  ;h  i�  ;h      H   ,  j�  ;h  j�  <0  kL  <0  kL  ;h  j�  ;h      H   ,  b�  ?P  b�  @  c|  @  c|  ?P  b�  ?P      H   ,  f�  =�  f�  >�  gd  >�  gd  =�  f�  =�      H   ,  e�  @�  e�  A�  f�  A�  f�  @�  e�  @�      H   ,  f�  ;h  f�  <0  gd  <0  gd  ;h  f�  ;h      H   ,  gd  =�  gd  >�  h,  >�  h,  =�  gd  =�      H   ,  c|  =�  c|  >�  dD  >�  dD  =�  c|  =�      H   ,  dD  <0  dD  <�  e  <�  e  <0  dD  <0      H   ,  gd  >�  gd  ?P  h,  ?P  h,  >�  gd  >�      H   ,  e�  <�  e�  =�  f�  =�  f�  <�  e�  <�      H   ,  dD  @�  dD  A�  e  A�  e  @�  dD  @�      H   ,  c|  <�  c|  =�  dD  =�  dD  <�  c|  <�      H   ,  c|  ?P  c|  @  dD  @  dD  ?P  c|  ?P      H   ,  dD  @  dD  @�  e  @�  e  @  dD  @      H   ,  e  <0  e  <�  e�  <�  e�  <0  e  <0      H   ,  gd  <�  gd  =�  h,  =�  h,  <�  gd  <�      H   ,  e  ?P  e  @  e�  @  e�  ?P  e  ?P      H   ,  e  ;h  e  <0  e�  <0  e�  ;h  e  ;h      H   ,  c|  <0  c|  <�  dD  <�  dD  <0  c|  <0      H   ,  dD  <�  dD  =�  e  =�  e  <�  dD  <�      H   ,  e  @  e  @�  e�  @�  e�  @  e  @      H   ,  b�  @�  b�  A�  c|  A�  c|  @�  b�  @�      H   ,  dD  ?P  dD  @  e  @  e  ?P  dD  ?P      H   ,  e�  @  e�  @�  f�  @�  f�  @  e�  @      H   ,  e�  =�  e�  >�  f�  >�  f�  =�  e�  =�      H   ,  b�  >�  b�  ?P  c|  ?P  c|  >�  b�  >�      H   ,  gd  <0  gd  <�  h,  <�  h,  <0  gd  <0      H   ,  e  <�  e  =�  e�  =�  e�  <�  e  <�      H   ,  f�  <�  f�  =�  gd  =�  gd  <�  f�  <�      H   ,  e�  ;h  e�  <0  f�  <0  f�  ;h  e�  ;h      H   ,  b�  =�  b�  >�  c|  >�  c|  =�  b�  =�      H   ,  e�  ?P  e�  @  f�  @  f�  ?P  e�  ?P      H   ,  dD  >�  dD  ?P  e  ?P  e  >�  dD  >�      H   ,  h,  =�  h,  >�  h�  >�  h�  =�  h,  =�      H   ,  gd  ;h  gd  <0  h,  <0  h,  ;h  gd  ;h      H   ,  f�  @  f�  @�  gd  @�  gd  @  f�  @      H   ,  e  @�  e  A�  e�  A�  e�  @�  e  @�      H   ,  e  =�  e  >�  e�  >�  e�  =�  e  =�      H   ,  h,  <�  h,  =�  h�  =�  h�  <�  h,  <�      H   ,  dD  =�  dD  >�  e  >�  e  =�  dD  =�      H   ,  e  >�  e  ?P  e�  ?P  e�  >�  e  >�      H   ,  c|  @�  c|  A�  dD  A�  dD  @�  c|  @�      H   ,  h,  <0  h,  <�  h�  <�  h�  <0  h,  <0      H   ,  c|  @  c|  @�  dD  @�  dD  @  c|  @      H   ,  f�  >�  f�  ?P  gd  ?P  gd  >�  f�  >�      H   ,  f�  ?P  f�  @  gd  @  gd  ?P  f�  ?P      H   ,  dD  ;h  dD  <0  e  <0  e  ;h  dD  ;h      H   ,  f�  <0  f�  <�  gd  <�  gd  <0  f�  <0      H   ,  h,  ;h  h,  <0  h�  <0  h�  ;h  h,  ;h      H   ,  b�  @  b�  @�  c|  @�  c|  @  b�  @      H   ,  e�  >�  e�  ?P  f�  ?P  f�  >�  e�  >�      H   ,  e�  <0  e�  <�  f�  <�  f�  <0  e�  <0      H   ,  c|  >�  c|  ?P  dD  ?P  dD  >�  c|  >�      H   ,  f�  9  f�  9�  gd  9�  gd  9  f�  9      H   ,  gd  9  gd  9�  h,  9�  h,  9  gd  9      H   ,  f�  9�  f�  :�  gd  :�  gd  9�  f�  9�      H   ,  e�  9�  e�  :�  f�  :�  f�  9�  e�  9�      H   ,  gd  8H  gd  9  h,  9  h,  8H  gd  8H      H   ,  h,  9  h,  9�  h�  9�  h�  9  h,  9      H   ,  h,  9�  h,  :�  h�  :�  h�  9�  h,  9�      H   ,  gd  9�  gd  :�  h,  :�  h,  9�  gd  9�      H   ,  h,  8H  h,  9  h�  9  h�  8H  h,  8H      H   ,  i�  9�  i�  :�  j�  :�  j�  9�  i�  9�      H   ,  o4  6�  o4  7�  o�  7�  o�  6�  o4  6�      H   ,  kL  9�  kL  :�  l  :�  l  9�  kL  9�      H   ,  nl  9  nl  9�  o4  9�  o4  9  nl  9      H   ,  l�  5(  l�  5�  m�  5�  m�  5(  l�  5(      H   ,  l  9  l  9�  l�  9�  l�  9  l  9      H   ,  m�  6�  m�  7�  nl  7�  nl  6�  m�  6�      H   ,  o4  8H  o4  9  o�  9  o�  8H  o4  8H      H   ,  j�  7�  j�  8H  kL  8H  kL  7�  j�  7�      H   ,  kL  7�  kL  8H  l  8H  l  7�  kL  7�      H   ,  kL  8H  kL  9  l  9  l  8H  kL  8H      H   ,  l�  6�  l�  7�  m�  7�  m�  6�  l�  6�      H   ,  i�  8H  i�  9  j�  9  j�  8H  i�  8H      H   ,  l  7�  l  8H  l�  8H  l�  7�  l  7�      H   ,  i�  9  i�  9�  j�  9�  j�  9  i�  9      H   ,  o4  7�  o4  8H  o�  8H  o�  7�  o4  7�      H   ,  l�  9�  l�  :�  m�  :�  m�  9�  l�  9�      H   ,  kL  6�  kL  7�  l  7�  l  6�  kL  6�      H   ,  j�  6�  j�  7�  kL  7�  kL  6�  j�  6�      H   ,  l  8H  l  9  l�  9  l�  8H  l  8H      H   ,  j�  9  j�  9�  kL  9�  kL  9  j�  9      H   ,  m�  5�  m�  6�  nl  6�  nl  5�  m�  5�      H   ,  m�  9�  m�  :�  nl  :�  nl  9�  m�  9�      H   ,  l  5�  l  6�  l�  6�  l�  5�  l  5�      H   ,  i�  7�  i�  8H  j�  8H  j�  7�  i�  7�      H   ,  nl  8H  nl  9  o4  9  o4  8H  nl  8H      H   ,  nl  9�  nl  :�  o4  :�  o4  9�  nl  9�      H   ,  nl  5�  nl  6�  o4  6�  o4  5�  nl  5�      H   ,  kL  5�  kL  6�  l  6�  l  5�  kL  5�      H   ,  o4  9  o4  9�  o�  9�  o�  9  o4  9      H   ,  l�  9  l�  9�  m�  9�  m�  9  l�  9      H   ,  j�  9�  j�  :�  kL  :�  kL  9�  j�  9�      H   ,  l�  5�  l�  6�  m�  6�  m�  5�  l�  5�      H   ,  nl  6�  nl  7�  o4  7�  o4  6�  nl  6�      H   ,  m�  7�  m�  8H  nl  8H  nl  7�  m�  7�      H   ,  m�  9  m�  9�  nl  9�  nl  9  m�  9      H   ,  nl  5(  nl  5�  o4  5�  o4  5(  nl  5(      H   ,  kL  9  kL  9�  l  9�  l  9  kL  9      H   ,  i�  6�  i�  7�  j�  7�  j�  6�  i�  6�      H   ,  j�  8H  j�  9  kL  9  kL  8H  j�  8H      H   ,  m�  8H  m�  9  nl  9  nl  8H  m�  8H      H   ,  o4  4`  o4  5(  o�  5(  o�  4`  o4  4`      H   ,  m�  5(  m�  5�  nl  5�  nl  5(  m�  5(      H   ,  l  6�  l  7�  l�  7�  l�  6�  l  6�      H   ,  l�  7�  l�  8H  m�  8H  m�  7�  l�  7�      H   ,  o4  5(  o4  5�  o�  5�  o�  5(  o4  5(      H   ,  nl  7�  nl  8H  o4  8H  o4  7�  nl  7�      H   ,  l  9�  l  :�  l�  :�  l�  9�  l  9�      H   ,  o4  5�  o4  6�  o�  6�  o�  5�  o4  5�      H   ,  l�  8H  l�  9  m�  9  m�  8H  l�  8H      H   ,  w�  2�  w�  3�  x�  3�  x�  2�  w�  2�      H   ,  y\  2  y\  2�  z$  2�  z$  2  y\  2      H   ,  ut  2�  ut  3�  v<  3�  v<  2�  ut  2�      H   ,  w  2�  w  3�  w�  3�  w�  2�  w  2�      H   ,  ||  2�  ||  3�  }D  3�  }D  2�  ||  2�      H   ,  s  2�  s  3�  s�  3�  s�  2�  s  2�      H   ,  z$  2  z$  2�  z�  2�  z�  2  z$  2      H   ,  }D  2  }D  2�  ~  2�  ~  2  }D  2      H   ,  s�  2�  s�  3�  t�  3�  t�  2�  s�  2�      H   ,  v<  2�  v<  3�  w  3�  w  2�  v<  2�      H   ,  x�  2�  x�  3�  y\  3�  y\  2�  x�  2�      H   ,  x�  1@  x�  2  y\  2  y\  1@  x�  1@      H   ,  y\  1@  y\  2  z$  2  z$  1@  y\  1@      H   ,  ut  2  ut  2�  v<  2�  v<  2  ut  2      H   ,  }D  0x  }D  1@  ~  1@  ~  0x  }D  0x      H   ,  z$  2�  z$  3�  z�  3�  z�  2�  z$  2�      H   ,  ||  2  ||  2�  }D  2�  }D  2  ||  2      H   ,  w  2  w  2�  w�  2�  w�  2  w  2      H   ,  }D  1@  }D  2  ~  2  ~  1@  }D  1@      H   ,  {�  0x  {�  1@  ||  1@  ||  0x  {�  0x      H   ,  x�  2  x�  2�  y\  2�  y\  2  x�  2      H   ,  y\  2�  y\  3�  z$  3�  z$  2�  y\  2�      H   ,  z$  1@  z$  2  z�  2  z�  1@  z$  1@      H   ,  {�  2�  {�  3�  ||  3�  ||  2�  {�  2�      H   ,  {�  1@  {�  2  ||  2  ||  1@  {�  1@      H   ,  }D  2�  }D  3�  ~  3�  ~  2�  }D  2�      H   ,  v<  2  v<  2�  w  2�  w  2  v<  2      H   ,  {�  2  {�  2�  ||  2�  ||  2  {�  2      H   ,  z�  2�  z�  3�  {�  3�  {�  2�  z�  2�      H   ,  z�  1@  z�  2  {�  2  {�  1@  z�  1@      H   ,  t�  2�  t�  3�  ut  3�  ut  2�  t�  2�      H   ,  w�  2  w�  2�  x�  2�  x�  2  w�  2      H   ,  ||  1@  ||  2  }D  2  }D  1@  ||  1@      H   ,  z�  2  z�  2�  {�  2�  {�  2  z�  2      H   ,  ||  0x  ||  1@  }D  1@  }D  0x  ||  0x      H   ,  }D  #�  }D  $�  ~  $�  ~  #�  }D  #�      H   ,  }D  @  }D    ~    ~  @  }D  @      H   ,  ||  �  ||  �  }D  �  }D  �  ||  �      H   ,  ||  x  ||  @  }D  @  }D  x  ||  x      H   ,  ||  �  ||  p  }D  p  }D  �  ||  �      H   ,  ||  (  ||  �  }D  �  }D  (  ||  (      H   ,  ||  H  ||     }D     }D  H  ||  H      H   ,  }D     }D  �  ~  �  ~     }D         H   ,  ||  �  ||  �  }D  �  }D  �  ||  �      H   ,  }D  �  }D  �  ~  �  ~  �  }D  �      H   ,  ||  `  ||  (  }D  (  }D  `  ||  `      H   ,  ||  �  ||  `  }D  `  }D  �  ||  �      H   ,  ||     ||  �  }D  �  }D     ||         H   ,  }D  !�  }D  "h  ~  "h  ~  !�  }D  !�      H   ,  }D  �  }D  x  ~  x  ~  �  }D  �      H   ,  }D  x  }D  @  ~  @  ~  x  }D  x      H   ,  }D  �  }D  H  ~  H  ~  �  }D  �      H   ,  {�  @  {�    ||    ||  @  {�  @      H   ,  {�     {�  �  ||  �  ||     {�         H   ,  }D    }D  �  ~  �  ~    }D        H   ,  }D     }D  �  ~  �  ~     }D         H   ,  ||  �  ||  X  }D  X  }D  �  ||  �      H   ,  }D  �  }D  �  ~  �  ~  �  }D  �      H   ,  }D  (  }D  �  ~  �  ~  (  }D  (      H   ,  }D  8  }D     ~     ~  8  }D  8      H   ,  }D  H  }D     ~     ~  H  }D  H      H   ,  }D  �  }D  X  ~  X  ~  �  }D  �      H   ,  }D  `  }D  (  ~  (  ~  `  }D  `      H   ,  ||  8  ||     }D     }D  8  ||  8      H   ,  }D  "h  }D  #0  ~  #0  ~  "h  }D  "h      H   ,  }D  p  }D  8  ~  8  ~  p  }D  p      H   ,  }D  X  }D     ~     ~  X  }D  X      H   ,  ||  @  ||    }D    }D  @  ||  @      H   ,  }D     }D   �  ~   �  ~     }D         H   ,  {�  x  {�  @  ||  @  ||  x  {�  x      H   ,  ||     ||  �  }D  �  }D     ||         H   ,  }D  �  }D  �  ~  �  ~  �  }D  �      H   ,  ||  �  ||  �  }D  �  }D  �  ||  �      H   ,  }D   �  }D  !�  ~  !�  ~   �  }D   �      H   ,  }D  �  }D  p  ~  p  ~  �  }D  �      H   ,  }D  �  }D  `  ~  `  ~  �  }D  �      H   ,  }D    }D  �  ~  �  ~    }D        H   ,  {�  �  {�  �  ||  �  ||  �  {�  �      H   ,  ||  �  ||  x  }D  x  }D  �  ||  �      H   ,  {�  �  {�  x  ||  x  ||  �  {�  �      H   ,  }D  �  }D  �  ~  �  ~  �  }D  �      H   ,  }D  �  }D  �  ~  �  ~  �  }D  �      H   ,  ||  p  ||  8  }D  8  }D  p  ||  p      H   ,  {�  �  {�  �  ||  �  ||  �  {�  �      H   ,  ||  �  ||  �  }D  �  }D  �  ||  �      H   ,  }D  �  }D  �  ~  �  ~  �  }D  �      H   ,  ||  �  ||  �  }D  �  }D  �  ||  �      H   ,  ||    ||  �  }D  �  }D    ||        H   ,  ||     ||   �  }D   �  }D     ||         H   ,  ||  �  ||  H  }D  H  }D  �  ||  �      H   ,  ||  X  ||     }D     }D  X  ||  X      H   ,  }D  #0  }D  #�  ~  #�  ~  #0  }D  #0      H   ,  {�    {�  �  ||  �  ||    {�        H   ,  {�  X  {�     ||     ||  X  {�  X      H   ,  �T  x  �T  @  �  @  �  x  �T  x      H   ,  ��  @  ��    �t    �t  @  ��  @      H   ,  �T  �  �T  x  �  x  �  �  �T  �      H   ,  ��  @  ��    ��    ��  @  ��  @      H   ,  �T  �  �T  �  �  �  �  �  �T  �      H   ,  �T     �T  �  �  �  �     �T         H   ,  �\  @  �\    �$    �$  @  �\  @      H   ,  �T  X  �T     �     �  X  �T  X      H   ,  �T  �  �T  X  �  X  �  �  �T  �      H   ,  �t  @  �t    �<    �<  @  �t  @      H   ,  �T  �  �T  �  �  �  �  �  �T  �      H   ,  �T     �T  �  �  �  �     �T         H   ,  �T  8  �T     �     �  8  �T  8      H   ,  ��  @  ��    ��    ��  @  ��  @      H   ,  �T  p  �T  8  �  8  �  p  �T  p      H   ,  �T  �  �T  p  �  p  �  �  �T  �      H   ,  ��  @  ��    �|    �|  @  ��  @      H   ,  �T  �  �T  �  �  �  �  �  �T  �      H   ,  ��  @  ��    ��    ��  @  ��  @      H   ,  �T    �T  �  �  �  �    �T        H   ,  �D  @  �D    �    �  @  �D  @      H   ,  �T  P  �T    �    �  P  �T  P      H   ,  ~�  @  ~�    �    �  @  ~�  @      H   ,  �T  �  �T  �  �  �  �  �  �T  �      H   ,  �  @  �    �d    �d  @  �  @      H   ,  �T  (  �T  �  �  �  �  (  �T  (      H   ,  �$  @  �$    ��    ��  @  �$  @      H   ,  �T  `  �T  (  �  (  �  `  �T  `      H   ,  �<  @  �<    �    �  @  �<  @      H   ,  ��  @  ��    ��    ��  @  ��  @      H   ,  �  @  �    ��    ��  @  �  @      H   ,  ��  @  ��    �\    �\  @  ��  @      H   ,  �4  @  �4    ��    ��  @  �4  @      H   ,  �T  �  �T  `  �  `  �  �  �T  �      H   ,  �  @  �    ��    ��  @  �  @      H   ,  �T  �  �T  �  �  �  �  �  �T  �      H   ,  ��  @  ��    �T    �T  @  ��  @      H   ,  ~  @  ~    ~�    ~�  @  ~  @      H   ,  �|  @  �|    �D    �D  @  �|  @      H   ,  �T    �T  �  �  �  �    �T        H   ,  �T  @  �T    �    �  @  �T  @      H   ,  ��  @  ��    ��    ��  @  ��  @      H   ,  ��  H  ��     �d     �d  H  ��  H      H   ,  �  H  �     ��     ��  H  �  H      H   ,  �\  �  �\  �  �$  �  �$  �  �\  �      H   ,  �\  �  �\  `  �$  `  �$  �  �\  �      H   ,  �\  �  �\  �  �$  �  �$  �  �\  �      H   ,  �D  H  �D     �     �  H  �D  H      H   ,  ��  H  ��     ��     ��  H  ��  H      H   ,  �\  `  �\  (  �$  (  �$  `  �\  `      H   ,  �\  (  �\  �  �$  �  �$  (  �\  (      H   ,  �\    �\  �  �$  �  �$    �\        H   ,  ��  !�  ��  "h  �d  "h  �d  !�  ��  !�      H   ,  ��  #�  ��  $�  �d  $�  �d  #�  ��  #�      H   ,  �|  %�  �|  &P  �D  &P  �D  %�  �|  %�      H   ,  �  $�  �  %�  ��  %�  ��  $�  �  $�      H   ,  �   �  �  !�  ��  !�  ��   �  �   �      H   ,  �|  $�  �|  %�  �D  %�  �D  $�  �|  $�      H   ,  ��  $�  ��  %�  �d  %�  �d  $�  ��  $�      H   ,  �D  #0  �D  #�  �  #�  �  #0  �D  #0      H   ,  �  #0  �  #�  ��  #�  ��  #0  �  #0      H   ,  ��     ��   �  �d   �  �d     ��         H   ,  ��  %�  ��  &P  ��  &P  ��  %�  ��  %�      H   ,  ��  #0  ��  #�  �d  #�  �d  #0  ��  #0      H   ,  �D  $�  �D  %�  �  %�  �  $�  �D  $�      H   ,  ��  $�  ��  %�  ��  %�  ��  $�  ��  $�      H   ,  �     �   �  ��   �  ��     �         H   ,  ��   �  ��  !�  �d  !�  �d   �  ��   �      H   ,  ��   �  ��  !�  ��  !�  ��   �  ��   �      H   ,  ��  "h  ��  #0  ��  #0  ��  "h  ��  "h      H   ,  �  "h  �  #0  ��  #0  ��  "h  �  "h      H   ,  ��  #�  ��  $�  ��  $�  ��  #�  ��  #�      H   ,  �  %�  �  &P  ��  &P  ��  %�  �  %�      H   ,  �  #�  �  $�  ��  $�  ��  #�  �  #�      H   ,  ��     ��   �  ��   �  ��     ��         H   ,  ��  %�  ��  &P  �|  &P  �|  %�  ��  %�      H   ,  �D  #�  �D  $�  �  $�  �  #�  �D  #�      H   ,  ��  #0  ��  #�  ��  #�  ��  #0  ��  #0      H   ,  ��  %�  ��  &P  �d  &P  �d  %�  ��  %�      H   ,  �D  %�  �D  &P  �  &P  �  %�  �D  %�      H   ,  ��  "h  ��  #0  �d  #0  �d  "h  ��  "h      H   ,  ��  !�  ��  "h  ��  "h  ��  !�  ��  !�      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  ��  `  ��  (  �t  (  �t  `  ��  `      H   ,  �  `  �  (  ��  (  ��  `  �  `      H   ,  ��    ��  �  �\  �  �\    ��        H   ,  �  (  �  �  ��  �  ��  (  �  (      H   ,  �<  �  �<  �  �  �  �  �  �<  �      H   ,  ��  �  ��  �  �t  �  �t  �  ��  �      H   ,  ��  �  ��  `  �\  `  �\  �  ��  �      H   ,  �  `  �  (  ��  (  ��  `  �  `      H   ,  �<    �<  �  �  �  �    �<        H   ,  �<  �  �<  �  �  �  �  �  �<  �      H   ,  ��  �  ��  `  ��  `  ��  �  ��  �      H   ,  ��  �  ��  `  �t  `  �t  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  �  ��  �  �\  �  �\  �  ��  �      H   ,  �  �  �  `  ��  `  ��  �  �  �      H   ,  �t  (  �t  �  �<  �  �<  (  �t  (      H   ,  �t    �t  �  �<  �  �<    �t        H   ,  ��  �  ��  �  �t  �  �t  �  ��  �      H   ,  �t  �  �t  `  �<  `  �<  �  �t  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��    ��  �  �t  �  �t    ��        H   ,  �    �  �  ��  �  ��    �        H   ,  ��  (  ��  �  �\  �  �\  (  ��  (      H   ,  �    �  �  ��  �  ��    �        H   ,  ��  `  ��  (  �\  (  �\  `  ��  `      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  `  ��  (  ��  (  ��  `  ��  `      H   ,  �<  (  �<  �  �  �  �  (  �<  (      H   ,  �<  �  �<  �  �  �  �  �  �<  �      H   ,  ��  (  ��  �  �t  �  �t  (  ��  (      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  `  ��  (  ��  (  ��  `  ��  `      H   ,  ��  (  ��  �  ��  �  ��  (  ��  (      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  ��  �  ��  `  ��  `  ��  �  ��  �      H   ,  �t  `  �t  (  �<  (  �<  `  �t  `      H   ,  �t  �  �t  �  �<  �  �<  �  �t  �      H   ,  �<  `  �<  (  �  (  �  `  �<  `      H   ,  ��  �  ��  �  �t  �  �t  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  �  ��  �  �\  �  �\  �  ��  �      H   ,  �t  �  �t  �  �<  �  �<  �  �t  �      H   ,  �  �  �  `  ��  `  ��  �  �  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �t  �  �t  �  �<  �  �<  �  �t  �      H   ,  �  (  �  �  ��  �  ��  (  �  (      H   ,  ��  (  ��  �  ��  �  ��  (  ��  (      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �<  �  �<  `  �  `  �  �  �<  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  H  ��  H  ��  �  ��  �      H   ,  �D  �  �D  �  �  �  �  �  �D  �      H   ,  �|  `  �|  (  �D  (  �D  `  �|  `      H   ,  �D  (  �D  �  �  �  �  (  �D  (      H   ,  �$  `  �$  (  ��  (  ��  `  �$  `      H   ,  ��  (  ��  �  ��  �  ��  (  ��  (      H   ,  ��  �  ��  �  �d  �  �d  �  ��  �      H   ,  �D    �D  �  �  �  �    �D        H   ,  �D  `  �D  (  �  (  �  `  �D  `      H   ,  ��  `  ��  (  �|  (  �|  `  ��  `      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �|  �  �|  `  �D  `  �D  �  �|  �      H   ,  �$  �  �$  `  ��  `  ��  �  �$  �      H   ,  �D  �  �D  `  �  `  �  �  �D  �      H   ,  ��  (  ��  �  �|  �  �|  (  ��  (      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �|  �  �|  �  �D  �  �D  �  �|  �      H   ,  ��  �  ��  H  �d  H  �d  �  ��  �      H   ,  ��  (  ��  �  �d  �  �d  (  ��  (      H   ,  �$  �  �$  �  ��  �  ��  �  �$  �      H   ,  �|  �  �|  H  �D  H  �D  �  �|  �      H   ,  �|    �|  �  �D  �  �D    �|        H   ,  �  `  �  (  ��  (  ��  `  �  `      H   ,  ��  �  ��  �  �|  �  �|  �  ��  �      H   ,  �$  �  �$  �  ��  �  ��  �  �$  �      H   ,  ��  `  ��  (  �d  (  �d  `  ��  `      H   ,  �    �  �  ��  �  ��    �        H   ,  �D  �  �D  H  �  H  �  �  �D  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  (  ��  �  ��  �  ��  (  ��  (      H   ,  ��  �  ��  `  ��  `  ��  �  ��  �      H   ,  �$    �$  �  ��  �  ��    �$        H   ,  �|  �  �|  �  �D  �  �D  �  �|  �      H   ,  ��  �  ��  `  �|  `  �|  �  ��  �      H   ,  ��    ��  �  �|  �  �|    ��        H   ,  �D  �  �D  �  �  �  �  �  �D  �      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  ��  �  ��  `  ��  `  ��  �  ��  �      H   ,  ��  �  ��  �  �d  �  �d  �  ��  �      H   ,  ��  `  ��  (  ��  (  ��  `  ��  `      H   ,  �|  �  �|  �  �D  �  �D  �  �|  �      H   ,  �  �  �  `  ��  `  ��  �  �  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �$  (  �$  �  ��  �  ��  (  �$  (      H   ,  �  �  �  H  ��  H  ��  �  �  �      H   ,  ��  `  ��  (  ��  (  ��  `  ��  `      H   ,  �  (  �  �  ��  �  ��  (  �  (      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  �  ��  �  �|  �  �|  �  ��  �      H   ,  ��  �  ��  �  �|  �  �|  �  ��  �      H   ,  �|  (  �|  �  �D  �  �D  (  �|  (      H   ,  �D  �  �D  �  �  �  �  �  �D  �      H   ,  �     �   �  �d   �  �d     �         H   ,  �d   �  �d  !�  �,  !�  �,   �  �d   �      H   ,  ~  �  ~  �  ~�  �  ~�  �  ~  �      H   ,  ��  `  ��  (  �T  (  �T  `  ��  `      H   ,  �  (  �  �  �d  �  �d  (  �  (      H   ,  �d  �  �d  �  �,  �  �,  �  �d  �      H   ,  ~�  �  ~�  �  �  �  �  �  ~�  �      H   ,  �d  !�  �d  "h  �,  "h  �,  !�  �d  !�      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  �    �  �  �d  �  �d    �        H   ,  ��    ��  �  �T  �  �T    ��        H   ,  ~�  �  ~�  H  �  H  �  �  ~�  �      H   ,  �  #0  �  #�  �d  #�  �d  #0  �  #0      H   ,  ~  `  ~  (  ~�  (  ~�  `  ~  `      H   ,  �,  %�  �,  &P  ��  &P  ��  %�  �,  %�      H   ,  ~  #�  ~  $�  ~�  $�  ~�  #�  ~  #�      H   ,  �d  H  �d     �,     �,  H  �d  H      H   ,  �d  "h  �d  #0  �,  #0  �,  "h  �d  "h      H   ,  ~  !�  ~  "h  ~�  "h  ~�  !�  ~  !�      H   ,  ��  %�  ��  &P  ��  &P  ��  %�  ��  %�      H   ,  ~�  %�  ~�  &P  �  &P  �  %�  ~�  %�      H   ,  ~�   �  ~�  !�  �  !�  �   �  ~�   �      H   ,  ��  (  ��  �  �T  �  �T  (  ��  (      H   ,  ~    ~  �  ~�  �  ~�    ~        H   ,  �d  %�  �d  &P  �,  &P  �,  %�  �d  %�      H   ,  ~�     ~�   �  �   �  �     ~�         H   ,  ~  #0  ~  #�  ~�  #�  ~�  #0  ~  #0      H   ,  ��  $�  ��  %�  ��  %�  ��  $�  ��  $�      H   ,  ~   �  ~  !�  ~�  !�  ~�   �  ~   �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �d  (  �d  �  �,  �  �,  (  �d  (      H   ,  ~�  $�  ~�  %�  �  %�  �  $�  ~�  $�      H   ,  ��  #�  ��  $�  ��  $�  ��  #�  ��  #�      H   ,  �d  #0  �d  #�  �,  #�  �,  #0  �d  #0      H   ,  �  !�  �  "h  �d  "h  �d  !�  �  !�      H   ,  �,  #�  �,  $�  ��  $�  ��  #�  �,  #�      H   ,  �  $�  �  %�  �d  %�  �d  $�  �  $�      H   ,  ��  �  ��  `  �T  `  �T  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ~  �  ~  H  ~�  H  ~�  �  ~  �      H   ,  ~�  �  ~�  �  �  �  �  �  ~�  �      H   ,  �,   �  �,  !�  ��  !�  ��   �  �,   �      H   ,  ~  �  ~  �  ~�  �  ~�  �  ~  �      H   ,  ~�  #�  ~�  $�  �  $�  �  #�  ~�  #�      H   ,  ~�  `  ~�  (  �  (  �  `  ~�  `      H   ,  ~�  !�  ~�  "h  �  "h  �  !�  ~�  !�      H   ,  �d  $�  �d  %�  �,  %�  �,  $�  �d  $�      H   ,  �,  "h  �,  #0  ��  #0  ��  "h  �,  "h      H   ,  �d  �  �d  �  �,  �  �,  �  �d  �      H   ,  ~  (  ~  �  ~�  �  ~�  (  ~  (      H   ,  ~  �  ~  `  ~�  `  ~�  �  ~  �      H   ,  �d     �d   �  �,   �  �,     �d         H   ,  �   �  �  !�  �d  !�  �d   �  �   �      H   ,  ~�  (  ~�  �  �  �  �  (  ~�  (      H   ,  �d  `  �d  (  �,  (  �,  `  �d  `      H   ,  �  H  �     �d     �d  H  �  H      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  ~�  H  ~�     �     �  H  ~�  H      H   ,  ��  �  ��  `  ��  `  ��  �  ��  �      H   ,  �,  !�  �,  "h  ��  "h  ��  !�  �,  !�      H   ,  �  `  �  (  �d  (  �d  `  �  `      H   ,  ~�  #0  ~�  #�  �  #�  �  #0  ~�  #0      H   ,  ��  `  ��  (  ��  (  ��  `  ��  `      H   ,  �,  #0  �,  #�  ��  #�  ��  #0  �,  #0      H   ,  �,  $�  �,  %�  ��  %�  ��  $�  �,  $�      H   ,  �d  #�  �d  $�  �,  $�  �,  #�  �d  #�      H   ,  �  �  �  �  �d  �  �d  �  �  �      H   ,  ~  �  ~  �  ~�  �  ~�  �  ~  �      H   ,  ~     ~   �  ~�   �  ~�     ~         H   ,  �  %�  �  &P  �d  &P  �d  %�  �  %�      H   ,  ~  $�  ~  %�  ~�  %�  ~�  $�  ~  $�      H   ,  ~�  �  ~�  �  �  �  �  �  ~�  �      H   ,  �  �  �  �  �d  �  �d  �  �  �      H   ,  ~�  "h  ~�  #0  �  #0  �  "h  ~�  "h      H   ,  ��  �  ��  �  �T  �  �T  �  ��  �      H   ,  ~�    ~�  �  �  �  �    ~�        H   ,  ~�  �  ~�  `  �  `  �  �  ~�  �      H   ,  �  �  �  H  �d  H  �d  �  �  �      H   ,  �  �  �  �  �d  �  �d  �  �  �      H   ,  �d  �  �d  H  �,  H  �,  �  �d  �      H   ,  ~  %�  ~  &P  ~�  &P  ~�  %�  ~  %�      H   ,  ~  H  ~     ~�     ~�  H  ~  H      H   ,  �  #�  �  $�  �d  $�  �d  #�  �  #�      H   ,  �  "h  �  #0  �d  #0  �d  "h  �  "h      H   ,  ~  "h  ~  #0  ~�  #0  ~�  "h  ~  "h      H   ,  �  �  �  `  �d  `  �d  �  �  �      H   ,  �L    �L  �  �  �  �    �L        H   ,  �L  �  �L  �  �  �  �  �  �L  �      H   ,  �  8  �     �d     �d  8  �  8      H   ,  ��  8  ��     ��     ��  8  ��  8      H   ,  ~  8  ~     ~�     ~�  8  ~  8      H   ,  �L  �  �L  �  �  �  �  �  �L  �      H   ,  �L  
�  �L  �  �  �  �  
�  �L  
�      H   ,  �d  8  �d     �,     �,  8  �d  8      H   ,  �L  P  �L    �    �  P  �L  P      H   ,  ~�  8  ~�     �     �  8  ~�  8      H   ,  ��  8  ��     ��     ��  8  ��  8      H   ,  �L  �  �L  P  �  P  �  �  �L  �      H   ,  ��  8  ��     �T     �T  8  ��  8      H   ,  ��  �  ��  x  �T  x  �T  �  ��  �      H   ,  ��  �  ��  X  ��  X  ��  �  ��  �      H   ,  ��  �  ��  X  �T  X  �T  �  ��  �      H   ,  �4  �  �4  X  ��  X  ��  �  �4  �      H   ,  �4     �4  �  ��  �  ��     �4         H   ,  ��  �  ��  �  �T  �  �T  �  ��  �      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  �4  X  �4     ��     ��  X  �4  X      H   ,  ��  x  ��  @  ��  @  ��  x  ��  x      H   ,  ��  �  ��  x  ��  x  ��  �  ��  �      H   ,  �4  x  �4  @  ��  @  ��  x  �4  x      H   ,  �4     �4  �  ��  �  ��     �4         H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��  X  ��     ��     ��  X  ��  X      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �4  �  �4  x  ��  x  ��  �  �4  �      H   ,  ��  x  ��  @  ��  @  ��  x  ��  x      H   ,  ��  X  ��     ��     ��  X  ��  X      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  x  ��  @  �T  @  �T  x  ��  x      H   ,  �4  �  �4  �  ��  �  ��  �  �4  �      H   ,  ��  X  ��     �T     �T  X  ��  X      H   ,  ��  �  ��  �  �T  �  �T  �  ��  �      H   ,  �4  �  �4  �  ��  �  ��  �  �4  �      H   ,  ��     ��  �  �T  �  �T     ��         H   ,  ��     ��  �  �T  �  �T     ��         H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  x  ��  x  ��  �  ��  �      H   ,  ��  �  ��  X  ��  X  ��  �  ��  �      H   ,  �  �  �  �  �d  �  �d  �  �  �      H   ,  ~�  X  ~�     �     �  X  ~�  X      H   ,  ~  �  ~  X  ~�  X  ~�  �  ~  �      H   ,  �d  �  �d  �  �,  �  �,  �  �d  �      H   ,  �  x  �  @  �d  @  �d  x  �  x      H   ,  ~�  �  ~�  X  �  X  �  �  ~�  �      H   ,  ~�  �  ~�  �  �  �  �  �  ~�  �      H   ,  ~  �  ~  x  ~�  x  ~�  �  ~  �      H   ,  �  �  �  X  �d  X  �d  �  �  �      H   ,  ~     ~  �  ~�  �  ~�     ~         H   ,  ~     ~  �  ~�  �  ~�     ~         H   ,  ~  x  ~  @  ~�  @  ~�  x  ~  x      H   ,  �     �  �  �d  �  �d     �         H   ,  ~  �  ~  �  ~�  �  ~�  �  ~  �      H   ,  ~�  x  ~�  @  �  @  �  x  ~�  x      H   ,  ~�     ~�  �  �  �  �     ~�         H   ,  �  X  �     �d     �d  X  �  X      H   ,  ~�  �  ~�  �  �  �  �  �  ~�  �      H   ,  �d     �d  �  �,  �  �,     �d         H   ,  ~�  �  ~�  x  �  x  �  �  ~�  �      H   ,  ~  �  ~  �  ~�  �  ~�  �  ~  �      H   ,  ~�     ~�  �  �  �  �     ~�         H   ,  ~  X  ~     ~�     ~�  X  ~  X      H   ,  �  �  �  x  �d  x  �d  �  �  �      H   ,  �     �  �  �d  �  �d     �         H   ,  �  �  �  �  �d  �  �d  �  �  �      H   ,  �d    �d  �  �,  �  �,    �d        H   ,  ~  P  ~    ~�    ~�  P  ~  P      H   ,  �  
�  �  �  �d  �  �d  
�  �  
�      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  �,  �  �,  �  ��  �  ��  �  �,  �      H   ,  ~�  �  ~�  p  �  p  �  �  ~�  �      H   ,  �,    �,  �  ��  �  ��    �,        H   ,  �,  
�  �,  �  ��  �  ��  
�  �,  
�      H   ,  �d  �  �d  P  �,  P  �,  �  �d  �      H   ,  ��  P  ��    �L    �L  P  ��  P      H   ,  �d  p  �d  8  �,  8  �,  p  �d  p      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  ~�    ~�  �  �  �  �    ~�        H   ,  �  p  �  8  �d  8  �d  p  �  p      H   ,  ~  �  ~  �  ~�  �  ~�  �  ~  �      H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  ��    ��  �  �L  �  �L    ��        H   ,  ��  
�  ��  �  �L  �  �L  
�  ��  
�      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �  �  �  �  �d  �  �d  �  �  �      H   ,  ��  �  ��  P  ��  P  ��  �  ��  �      H   ,  �,  P  �,    ��    ��  P  �,  P      H   ,  ��  �  ��  �  �L  �  �L  �  ��  �      H   ,  �d  P  �d    �,    �,  P  �d  P      H   ,  ~�  �  ~�  �  �  �  �  �  ~�  �      H   ,  ~  �  ~  p  ~�  p  ~�  �  ~  �      H   ,  �  �  �  �  �d  �  �d  �  �  �      H   ,  �,  p  �,  8  ��  8  ��  p  �,  p      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  P  ��  P  ��  �  ��  �      H   ,  �  �  �  P  �d  P  �d  �  �  �      H   ,  ~  �  ~  P  ~�  P  ~�  �  ~  �      H   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      H   ,  �d  
�  �d  �  �,  �  �,  
�  �d  
�      H   ,  �d  �  �d  p  �,  p  �,  �  �d  �      H   ,  �  �  �  p  �d  p  �d  �  �  �      H   ,  ~�  p  ~�  8  �  8  �  p  ~�  p      H   ,  ��  �  ��  P  �L  P  �L  �  ��  �      H   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      H   ,  ~�  P  ~�    �    �  P  ~�  P      H   ,  ~    ~  �  ~�  �  ~�    ~        H   ,  �,  �  �,  P  ��  P  ��  �  �,  �      H   ,  �,  �  �,  �  ��  �  ��  �  �,  �      H   ,  ~�  �  ~�  P  �  P  �  �  ~�  �      H   ,  ~�  �  ~�  �  �  �  �  �  ~�  �      H   ,  �d  �  �d  �  �,  �  �,  �  �d  �      H   ,  �  P  �    �d    �d  P  �  P      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ~  p  ~  8  ~�  8  ~�  p  ~  p      H   ,  �,  �  �,  p  ��  p  ��  �  �,  �      H   ,  �    �  �  �d  �  �d    �        H   ,  �d  �  �d  �  �,  �  �,  �  �d  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  p  �l  p  �l  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  �  ��  P  �T  P  �T  �  ��  �      H   ,  ��  �  ��  �  �l  �  �l  �  ��  �      H   ,  �4    �4  �  ��  �  ��    �4        H   ,  �4  P  �4    ��    ��  P  �4  P      H   ,  �l  �  �l  �  �4  �  �4  �  �l  �      H   ,  ��  p  ��  8  �T  8  �T  p  ��  p      H   ,  �  �  �  P  ��  P  ��  �  �  �      H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  �  
�  �  �  ��  �  ��  
�  �  
�      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  �l  �  �l  �  �4  �  �4  �  �l  �      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  �l    �l  �  �4  �  �4    �l        H   ,  ��  �  ��  p  �T  p  �T  �  ��  �      H   ,  ��  �  ��  �  �T  �  �T  �  ��  �      H   ,  ��  
�  ��  �  �l  �  �l  
�  ��  
�      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  P  ��    �T    �T  P  ��  P      H   ,  �l  �  �l  P  �4  P  �4  �  �l  �      H   ,  ��  �  ��  P  ��  P  ��  �  ��  �      H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  �4  p  �4  8  ��  8  ��  p  �4  p      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  �l  P  �l    �4    �4  P  �l  P      H   ,  �    �  �  ��  �  ��    �        H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  �  �l  �  �l  �  ��  �      H   ,  �l  �  �l  p  �4  p  �4  �  �l  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �4  �  �4  p  ��  p  ��  �  �4  �      H   ,  �  P  �    ��    ��  P  �  P      H   ,  �4  �  �4  �  ��  �  ��  �  �4  �      H   ,  �l  
�  �l  �  �4  �  �4  
�  �l  
�      H   ,  �4  �  �4  �  ��  �  ��  �  �4  �      H   ,  ��    ��  �  �l  �  �l    ��        H   ,  ��    ��  �  ��  �  ��    ��        H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  
�  ��  �  ��  �  ��  
�  ��  
�      H   ,  ��  �  ��  P  ��  P  ��  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  �4  �  �4  P  ��  P  ��  �  �4  �      H   ,  ��    ��  �  �T  �  �T    ��        H   ,  ��  �  ��  P  �l  P  �l  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  P  ��  P  ��  �  ��  �      H   ,  ��  P  ��    �l    �l  P  ��  P      H   ,  �\  P  �\    �$    �$  P  �\  P      H   ,  ��  8  ��     ��     ��  8  ��  8      H   ,  �\  �  �\  �  �$  �  �$  �  �\  �      H   ,  �\  �  �\  �  �$  �  �$  �  �\  �      H   ,  �\  �  �\  x  �$  x  �$  �  �\  �      H   ,  �\  X  �\     �$     �$  X  �\  X      H   ,  �  8  �     ��     ��  8  �  8      H   ,  ��  8  ��     ��     ��  8  ��  8      H   ,  �\     �\  �  �$  �  �$     �\         H   ,  �$  8  �$     ��     ��  8  �$  8      H   ,  ��  8  ��     �\     �\  8  ��  8      H   ,  ��  8  ��     �t     �t  8  ��  8      H   ,  �\  �  �\  p  �$  p  �$  �  �\  �      H   ,  �\    �\  �  �$  �  �$    �\        H   ,  �<  8  �<     �     �  8  �<  8      H   ,  ��  8  ��     ��     ��  8  ��  8      H   ,  �\     �\  �  �$  �  �$     �\         H   ,  �\  �  �\  X  �$  X  �$  �  �\  �      H   ,  �|  8  �|     �D     �D  8  �|  8      H   ,  �\  �  �\  �  �$  �  �$  �  �\  �      H   ,  �\  8  �\     �$     �$  8  �\  8      H   ,  ��  8  ��     �|     �|  8  ��  8      H   ,  �  8  �     ��     ��  8  �  8      H   ,  �t  8  �t     �<     �<  8  �t  8      H   ,  �\  p  �\  8  �$  8  �$  p  �\  p      H   ,  �\  x  �\  @  �$  @  �$  x  �\  x      H   ,  �$     �$  �  ��  �  ��     �$         H   ,  �|     �|  �  �D  �  �D     �|         H   ,  �|  X  �|     �D     �D  X  �|  X      H   ,  �     �  �  ��  �  ��     �         H   ,  ��  �  ��  X  �|  X  �|  �  ��  �      H   ,  �|  �  �|  �  �D  �  �D  �  �|  �      H   ,  �$  X  �$     ��     ��  X  �$  X      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��  �  ��  x  �|  x  �|  �  ��  �      H   ,  �D  �  �D  X  �  X  �  �  �D  �      H   ,  ��     ��  �  �|  �  �|     ��         H   ,  ��  x  ��  @  �|  @  �|  x  ��  x      H   ,  ��  X  ��     ��     ��  X  ��  X      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��     ��  �  �|  �  �|     ��         H   ,  ��  �  ��  X  ��  X  ��  �  ��  �      H   ,  �|  �  �|  �  �D  �  �D  �  �|  �      H   ,  �$     �$  �  ��  �  ��     �$         H   ,  �$  �  �$  X  ��  X  ��  �  �$  �      H   ,  ��  �  ��  x  ��  x  ��  �  ��  �      H   ,  �D     �D  �  �  �  �     �D         H   ,  �$  x  �$  @  ��  @  ��  x  �$  x      H   ,  �|  x  �|  @  �D  @  �D  x  �|  x      H   ,  �D  �  �D  �  �  �  �  �  �D  �      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  �D  x  �D  @  �  @  �  x  �D  x      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �|     �|  �  �D  �  �D     �|         H   ,  �$  �  �$  x  ��  x  ��  �  �$  �      H   ,  �D     �D  �  �  �  �     �D         H   ,  ��  �  ��  �  �|  �  �|  �  ��  �      H   ,  ��  x  ��  @  ��  @  ��  x  ��  x      H   ,  �$  �  �$  �  ��  �  ��  �  �$  �      H   ,  �|  �  �|  x  �D  x  �D  �  �|  �      H   ,  �D  �  �D  �  �  �  �  �  �D  �      H   ,  ��  �  ��  �  �|  �  �|  �  ��  �      H   ,  �D  X  �D     �     �  X  �D  X      H   ,  �D  �  �D  x  �  x  �  �  �D  �      H   ,  �|  �  �|  X  �D  X  �D  �  �|  �      H   ,  ��  X  ��     �|     �|  X  ��  X      H   ,  �$  �  �$  �  ��  �  ��  �  �$  �      H   ,  �t  �  �t  X  �<  X  �<  �  �t  �      H   ,  �<  �  �<  x  �  x  �  �  �<  �      H   ,  ��  X  ��     �t     �t  X  ��  X      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  �  ��  X  �t  X  �t  �  ��  �      H   ,  �  �  �  x  ��  x  ��  �  �  �      H   ,  �<  X  �<     �     �  X  �<  X      H   ,  ��  �  ��  x  �t  x  �t  �  ��  �      H   ,  �<  �  �<  �  �  �  �  �  �<  �      H   ,  ��  X  ��     �\     �\  X  ��  X      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  �     �  �  ��  �  ��     �         H   ,  �  �  �  X  ��  X  ��  �  �  �      H   ,  �t     �t  �  �<  �  �<     �t         H   ,  ��  �  ��  �  �\  �  �\  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��     ��  �  �t  �  �t     ��         H   ,  ��  �  ��  x  ��  x  ��  �  ��  �      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��  �  ��  x  ��  x  ��  �  ��  �      H   ,  ��  �  ��  X  �\  X  �\  �  ��  �      H   ,  ��  �  ��  �  �t  �  �t  �  ��  �      H   ,  ��     ��  �  �\  �  �\     ��         H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �<  �  �<  X  �  X  �  �  �<  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �     �  �  ��  �  ��     �         H   ,  ��  �  ��  X  ��  X  ��  �  ��  �      H   ,  �     �  �  ��  �  ��     �         H   ,  �  �  �  X  ��  X  ��  �  �  �      H   ,  ��  X  ��     ��     ��  X  ��  X      H   ,  �t  �  �t  �  �<  �  �<  �  �t  �      H   ,  ��     ��  �  �\  �  �\     ��         H   ,  ��  �  ��  X  ��  X  ��  �  ��  �      H   ,  ��  x  ��  @  ��  @  ��  x  ��  x      H   ,  �  X  �     ��     ��  X  �  X      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  x  �\  x  �\  �  ��  �      H   ,  �  x  �  @  ��  @  ��  x  �  x      H   ,  ��  X  ��     ��     ��  X  ��  X      H   ,  ��  x  ��  @  �t  @  �t  x  ��  x      H   ,  ��  �  ��  �  �\  �  �\  �  ��  �      H   ,  �t  �  �t  x  �<  x  �<  �  �t  �      H   ,  �  �  �  x  ��  x  ��  �  �  �      H   ,  �t  x  �t  @  �<  @  �<  x  �t  x      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �  x  �  @  ��  @  ��  x  �  x      H   ,  �<     �<  �  �  �  �     �<         H   ,  �t  X  �t     �<     �<  X  �t  X      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �     �  �  ��  �  ��     �         H   ,  �<  �  �<  �  �  �  �  �  �<  �      H   ,  �<     �<  �  �  �  �     �<         H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��  x  ��  @  ��  @  ��  x  ��  x      H   ,  ��     ��  �  �t  �  �t     ��         H   ,  ��  �  ��  �  �t  �  �t  �  ��  �      H   ,  �t  �  �t  �  �<  �  �<  �  �t  �      H   ,  �  X  �     ��     ��  X  �  X      H   ,  ��  x  ��  @  �\  @  �\  x  ��  x      H   ,  �t     �t  �  �<  �  �<     �t         H   ,  �<  x  �<  @  �  @  �  x  �<  x      H   ,  �t    �t  �  �<  �  �<    �t        H   ,  ��  �  ��  �  �\  �  �\  �  ��  �      H   ,  �t  �  �t  �  �<  �  �<  �  �t  �      H   ,  �t  p  �t  8  �<  8  �<  p  �t  p      H   ,  ��  P  ��    �\    �\  P  ��  P      H   ,  �t  �  �t  p  �<  p  �<  �  �t  �      H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  �<  �  �<  p  �  p  �  �  �<  �      H   ,  �    �  �  ��  �  ��    �        H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �  P  �    ��    ��  P  �  P      H   ,  ��    ��  �  �t  �  �t    ��        H   ,  �  �  �  p  ��  p  ��  �  �  �      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �  p  �  8  ��  8  ��  p  �  p      H   ,  ��  p  ��  8  �t  8  �t  p  ��  p      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �<  P  �<    �    �  P  �<  P      H   ,  �<  p  �<  8  �  8  �  p  �<  p      H   ,  ��  P  ��    �t    �t  P  ��  P      H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  ��  �  ��  p  �\  p  �\  �  ��  �      H   ,  ��  �  ��  p  �t  p  �t  �  ��  �      H   ,  �  p  �  8  ��  8  ��  p  �  p      H   ,  �<    �<  �  �  �  �    �<        H   ,  �  �  �  p  ��  p  ��  �  �  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��    ��  �  �\  �  �\    ��        H   ,  �    �  �  ��  �  ��    �        H   ,  ��    ��  �  ��  �  ��    ��        H   ,  �<  �  �<  �  �  �  �  �  �<  �      H   ,  ��  �  ��  �  �t  �  �t  �  ��  �      H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  �t  P  �t    �<    �<  P  �t  P      H   ,  ��  p  ��  8  �\  8  �\  p  ��  p      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  �$  �  �$  p  ��  p  ��  �  �$  �      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  ��  p  ��  8  �|  8  �|  p  ��  p      H   ,  �|  p  �|  8  �D  8  �D  p  �|  p      H   ,  �$  �  �$  �  ��  �  ��  �  �$  �      H   ,  �$    �$  �  ��  �  ��    �$        H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �$  p  �$  8  ��  8  ��  p  �$  p      H   ,  ��  �  ��  p  �|  p  �|  �  ��  �      H   ,  �  6�  �  7�  ��  7�  ��  6�  �  6�      H   ,  �  3�  �  4`  ��  4`  ��  3�  �  3�      H   ,  �  5�  �  6�  ��  6�  ��  5�  �  5�      H   ,  �  5(  �  5�  ��  5�  ��  5(  �  5(      H   ,  �  4`  �  5(  ��  5(  ��  4`  �  4`      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  �l  3�  �l  4`  �4  4`  �4  3�  �l  3�      H   ,  �<  3�  �<  4`  �  4`  �  3�  �<  3�      H   ,  �4  3�  �4  4`  ��  4`  ��  3�  �4  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  �T  3�  �T  4`  �  4`  �  3�  �T  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  �L  3�  �L  4`  �  4`  �  3�  �L  3�      H   ,  ��  3�  ��  4`  �L  4`  �L  3�  ��  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  ��  3�  ��  4`  �l  4`  �l  3�  ��  3�      H   ,  �t  3�  �t  4`  �<  4`  �<  3�  �t  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  �  @�  �  A�  ��  A�  ��  @�  �  @�      H   ,  �  @  �  @�  ��  @�  ��  @  �  @      H   ,  �  3�  �  4`  ��  4`  ��  3�  �  3�      H   ,  ��  3�  ��  4`  �T  4`  �T  3�  ��  3�      H   ,  �  8H  �  9  ��  9  ��  8H  �  8H      H   ,  ��  3�  ��  4`  �t  4`  �t  3�  ��  3�      H   ,  �  7�  �  8H  ��  8H  ��  7�  �  7�      H   ,  ��  :�  ��  ;h  ƴ  ;h  ƴ  :�  ��  :�      H   ,  �d  :�  �d  ;h  �,  ;h  �,  :�  �d  :�      H   ,  ��  :�  ��  ;h  ͼ  ;h  ͼ  :�  ��  :�      H   ,  �  <�  �  =�  ��  =�  ��  <�  �  <�      H   ,  �  <0  �  <�  ��  <�  ��  <0  �  <0      H   ,  �  ;h  �  <0  ��  <0  ��  ;h  �  ;h      H   ,  �  :�  �  ;h  ��  ;h  ��  :�  �  :�      H   ,  ʜ  :�  ʜ  ;h  �d  ;h  �d  :�  ʜ  :�      H   ,  �  9�  �  :�  ��  :�  ��  9�  �  9�      H   ,  �D  :�  �D  ;h  �  ;h  �  :�  �D  :�      H   ,  �  9  �  9�  ��  9�  ��  9  �  9      H   ,  ͼ  :�  ͼ  ;h  ΄  ;h  ΄  :�  ͼ  :�      H   ,  ��  :�  ��  ;h  ʜ  ;h  ʜ  :�  ��  :�      H   ,  ƴ  :�  ƴ  ;h  �|  ;h  �|  :�  ƴ  :�      H   ,  �  8H  �  9  ��  9  ��  8H  �  8H      H   ,  �|  :�  �|  ;h  �D  ;h  �D  :�  �|  :�      H   ,  �  7�  �  8H  ��  8H  ��  7�  �  7�      H   ,  �,  :�  �,  ;h  ��  ;h  ��  :�  �,  :�      H   ,  ��  <�  ��  =�  ͼ  =�  ͼ  <�  ��  <�      H   ,  ΄  >�  ΄  ?P  �L  ?P  �L  >�  ΄  >�      H   ,  ��  <0  ��  <�  ͼ  <�  ͼ  <0  ��  <0      H   ,  ��  @�  ��  A�  ͼ  A�  ͼ  @�  ��  @�      H   ,  ��  ;h  ��  <0  ͼ  <0  ͼ  ;h  ��  ;h      H   ,  �d  =�  �d  >�  �,  >�  �,  =�  �d  =�      H   ,  ΄  =�  ΄  >�  �L  >�  �L  =�  ΄  =�      H   ,  ΄  <�  ΄  =�  �L  =�  �L  <�  ΄  <�      H   ,  �L  @�  �L  A�  �  A�  �  @�  �L  @�      H   ,  ʜ  >�  ʜ  ?P  �d  ?P  �d  >�  ʜ  >�      H   ,  ΄  @  ΄  @�  �L  @�  �L  @  ΄  @      H   ,  ʜ  =�  ʜ  >�  �d  >�  �d  =�  ʜ  =�      H   ,  ��  @  ��  @�  ͼ  @�  ͼ  @  ��  @      H   ,  ʜ  <�  ʜ  =�  �d  =�  �d  <�  ʜ  <�      H   ,  ΄  <0  ΄  <�  �L  <�  �L  <0  ΄  <0      H   ,  ʜ  <0  ʜ  <�  �d  <�  �d  <0  ʜ  <0      H   ,  �L  @  �L  @�  �  @�  �  @  �L  @      H   ,  ͼ  @�  ͼ  A�  ΄  A�  ΄  @�  ͼ  @�      H   ,  ʜ  ;h  ʜ  <0  �d  <0  �d  ;h  ʜ  ;h      H   ,  ��  =�  ��  >�  ʜ  >�  ʜ  =�  ��  =�      H   ,  ͼ  @  ͼ  @�  ΄  @�  ΄  @  ͼ  @      H   ,  �d  <�  �d  =�  �,  =�  �,  <�  �d  <�      H   ,  �L  ?P  �L  @  �  @  �  ?P  �L  ?P      H   ,  ͼ  ?P  ͼ  @  ΄  @  ΄  ?P  ͼ  ?P      H   ,  ��  <�  ��  =�  ʜ  =�  ʜ  <�  ��  <�      H   ,  ͼ  >�  ͼ  ?P  ΄  ?P  ΄  >�  ͼ  >�      H   ,  ��  ?P  ��  @  ͼ  @  ͼ  ?P  ��  ?P      H   ,  �L  >�  �L  ?P  �  ?P  �  >�  �L  >�      H   ,  ͼ  =�  ͼ  >�  ΄  >�  ΄  =�  ͼ  =�      H   ,  �,  @�  �,  A�  ��  A�  ��  @�  �,  @�      H   ,  ��  <0  ��  <�  ʜ  <�  ʜ  <0  ��  <0      H   ,  ͼ  <�  ͼ  =�  ΄  =�  ΄  <�  ͼ  <�      H   ,  �,  @  �,  @�  ��  @�  ��  @  �,  @      H   ,  ͼ  <0  ͼ  <�  ΄  <�  ΄  <0  ͼ  <0      H   ,  ��  ;h  ��  <0  ʜ  <0  ʜ  ;h  ��  ;h      H   ,  �,  ?P  �,  @  ��  @  ��  ?P  �,  ?P      H   ,  ��  >�  ��  ?P  ͼ  ?P  ͼ  >�  ��  >�      H   ,  ͼ  ;h  ͼ  <0  ΄  <0  ΄  ;h  ͼ  ;h      H   ,  �,  >�  �,  ?P  ��  ?P  ��  >�  �,  >�      H   ,  ΄  ?P  ΄  @  �L  @  �L  ?P  ΄  ?P      H   ,  �d  <0  �d  <�  �,  <�  �,  <0  �d  <0      H   ,  �,  =�  �,  >�  ��  >�  ��  =�  �,  =�      H   ,  �L  =�  �L  >�  �  >�  �  =�  �L  =�      H   ,  ��  =�  ��  >�  ͼ  >�  ͼ  =�  ��  =�      H   ,  �,  <�  �,  =�  ��  =�  ��  <�  �,  <�      H   ,  �d  ?P  �d  @  �,  @  �,  ?P  �d  ?P      H   ,  �,  <0  �,  <�  ��  <�  ��  <0  �,  <0      H   ,  �L  <�  �L  =�  �  =�  �  <�  �L  <�      H   ,  �d  ;h  �d  <0  �,  <0  �,  ;h  �d  ;h      H   ,  �,  ;h  �,  <0  ��  <0  ��  ;h  �,  ;h      H   ,  �d  >�  �d  ?P  �,  ?P  �,  >�  �d  >�      H   ,  ΄  @�  ΄  A�  �L  A�  �L  @�  ΄  @�      H   ,  ƴ  ;h  ƴ  <0  �|  <0  �|  ;h  ƴ  ;h      H   ,  Ô  @�  Ô  A�  �\  A�  �\  @�  Ô  @�      H   ,  �|  ;h  �|  <0  �D  <0  �D  ;h  �|  ;h      H   ,  ��  @  ��  @�  ƴ  @�  ƴ  @  ��  @      H   ,  ��  @�  ��  A�  Ô  A�  Ô  @�  ��  @�      H   ,  �\  @  �\  @�  �$  @�  �$  @  �\  @      H   ,  �D  ;h  �D  <0  �  <0  �  ;h  �D  ;h      H   ,  �$  @�  �$  A�  ��  A�  ��  @�  �$  @�      H   ,  �D  <0  �D  <�  �  <�  �  <0  �D  <0      H   ,  ��  @�  ��  A�  ƴ  A�  ƴ  @�  ��  @�      H   ,  Ô  @  Ô  @�  �\  @�  �\  @  Ô  @      H   ,  �\  @�  �\  A�  �$  A�  �$  @�  �\  @�      H   ,  ƴ  @�  ƴ  A�  �|  A�  �|  @�  ƴ  @�      H   ,  �$  @  �$  @�  ��  @�  ��  @  �$  @      H   ,  ��  @  ��  @�  Ô  @�  Ô  @  ��  @      H   ,  �|  @�  �|  A�  �D  A�  �D  @�  �|  @�      H   ,  �|  9�  �|  :�  �D  :�  �D  9�  �|  9�      H   ,  Ô  7�  Ô  8H  �\  8H  �\  7�  Ô  7�      H   ,  �\  9  �\  9�  �$  9�  �$  9  �\  9      H   ,  �|  8H  �|  9  �D  9  �D  8H  �|  8H      H   ,  �$  9�  �$  :�  ��  :�  ��  9�  �$  9�      H   ,  Ô  8H  Ô  9  �\  9  �\  8H  Ô  8H      H   ,  �\  5(  �\  5�  �$  5�  �$  5(  �\  5(      H   ,  �\  8H  �\  9  �$  9  �$  8H  �\  8H      H   ,  �$  9  �$  9�  ��  9�  ��  9  �$  9      H   ,  �D  8H  �D  9  �  9  �  8H  �D  8H      H   ,  �D  7�  �D  8H  �  8H  �  7�  �D  7�      H   ,  �\  5�  �\  6�  �$  6�  �$  5�  �\  5�      H   ,  ��  9�  ��  :�  ƴ  :�  ƴ  9�  ��  9�      H   ,  ��  8H  ��  9  Ô  9  Ô  8H  ��  8H      H   ,  �|  6�  �|  7�  �D  7�  �D  6�  �|  6�      H   ,  �$  8H  �$  9  ��  9  ��  8H  �$  8H      H   ,  �|  9  �|  9�  �D  9�  �D  9  �|  9      H   ,  Ô  6�  Ô  7�  �\  7�  �\  6�  Ô  6�      H   ,  ��  9  ��  9�  Ô  9�  Ô  9  ��  9      H   ,  �$  7�  �$  8H  ��  8H  ��  7�  �$  7�      H   ,  ��  6�  ��  7�  Ô  7�  Ô  6�  ��  6�      H   ,  ��  9  ��  9�  ƴ  9�  ƴ  9  ��  9      H   ,  �|  7�  �|  8H  �D  8H  �D  7�  �|  7�      H   ,  �D  9�  �D  :�  �  :�  �  9�  �D  9�      H   ,  ��  8H  ��  9  ƴ  9  ƴ  8H  ��  8H      H   ,  Ô  9  Ô  9�  �\  9�  �\  9  Ô  9      H   ,  �$  6�  �$  7�  ��  7�  ��  6�  �$  6�      H   ,  Ô  5�  Ô  6�  �\  6�  �\  5�  Ô  5�      H   ,  ��  7�  ��  8H  ƴ  8H  ƴ  7�  ��  7�      H   ,  ƴ  9�  ƴ  :�  �|  :�  �|  9�  ƴ  9�      H   ,  �\  7�  �\  8H  �$  8H  �$  7�  �\  7�      H   ,  ��  5�  ��  6�  Ô  6�  Ô  5�  ��  5�      H   ,  �$  5�  �$  6�  ��  6�  ��  5�  �$  5�      H   ,  ƴ  9  ƴ  9�  �|  9�  �|  9  ƴ  9      H   ,  ƴ  8H  ƴ  9  �|  9  �|  8H  ƴ  8H      H   ,  �D  6�  �D  7�  �  7�  �  6�  �D  6�      H   ,  �$  5(  �$  5�  ��  5�  ��  5(  �$  5(      H   ,  ��  6�  ��  7�  ƴ  7�  ƴ  6�  ��  6�      H   ,  Ô  5(  Ô  5�  �\  5�  �\  5(  Ô  5(      H   ,  ƴ  7�  ƴ  8H  �|  8H  �|  7�  ƴ  7�      H   ,  �\  6�  �\  7�  �$  7�  �$  6�  �\  6�      H   ,  ��  5�  ��  6�  ƴ  6�  ƴ  5�  ��  5�      H   ,  ��  5(  ��  5�  Ô  5�  Ô  5(  ��  5(      H   ,  ƴ  6�  ƴ  7�  �|  7�  �|  6�  ƴ  6�      H   ,  �\  9�  �\  :�  �$  :�  �$  9�  �\  9�      H   ,  ƴ  5�  ƴ  6�  �|  6�  �|  5�  ƴ  5�      H   ,  Ô  4`  Ô  5(  �\  5(  �\  4`  Ô  4`      H   ,  ��  7�  ��  8H  Ô  8H  Ô  7�  ��  7�      H   ,  �D  9  �D  9�  �  9�  �  9  �D  9      H   ,  ��  4`  ��  5(  Ô  5(  Ô  4`  ��  4`      H   ,  ʜ  9�  ʜ  :�  �d  :�  �d  9�  ʜ  9�      H   ,  ʜ  8H  ʜ  9  �d  9  �d  8H  ʜ  8H      H   ,  �d  9  �d  9�  �,  9�  �,  9  �d  9      H   ,  ��  9  ��  9�  ʜ  9�  ʜ  9  ��  9      H   ,  ʜ  9  ʜ  9�  �d  9�  �d  9  ʜ  9      H   ,  ��  9�  ��  :�  ͼ  :�  ͼ  9�  ��  9�      H   ,  ��  7�  ��  8H  ʜ  8H  ʜ  7�  ��  7�      H   ,  �,  9�  �,  :�  ��  :�  ��  9�  �,  9�      H   ,  �d  9�  �d  :�  �,  :�  �,  9�  �d  9�      H   ,  ��  8H  ��  9  ʜ  9  ʜ  8H  ��  8H      H   ,  ��  9�  ��  :�  ʜ  :�  ʜ  9�  ��  9�      H   ,  �T  5�  �T  6�  �  6�  �  5�  �T  5�      H   ,  ��  6�  ��  7�  �T  7�  �T  6�  ��  6�      H   ,  �l  5(  �l  5�  �4  5�  �4  5(  �l  5(      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  �<  5(  �<  5�  �  5�  �  5(  �<  5(      H   ,  �l  5�  �l  6�  �4  6�  �4  5�  �l  5�      H   ,  ��  6�  ��  7�  ��  7�  ��  6�  ��  6�      H   ,  �4  4`  �4  5(  ��  5(  ��  4`  �4  4`      H   ,  ��  5�  ��  6�  �l  6�  �l  5�  ��  5�      H   ,  �  5(  �  5�  ��  5�  ��  5(  �  5(      H   ,  ��  5�  ��  6�  �T  6�  �T  5�  ��  5�      H   ,  �T  5(  �T  5�  �  5�  �  5(  �T  5(      H   ,  �<  7�  �<  8H  �  8H  �  7�  �<  7�      H   ,  �4  5(  �4  5�  ��  5�  ��  5(  �4  5(      H   ,  �L  4`  �L  5(  �  5(  �  4`  �L  4`      H   ,  �<  @�  �<  A�  �  A�  �  @�  �<  @�      H   ,  ��  4`  ��  5(  �l  5(  �l  4`  ��  4`      H   ,  ��  5�  ��  6�  ��  6�  ��  5�  ��  5�      H   ,  �  4`  �  5(  ��  5(  ��  4`  �  4`      H   ,  ��  5(  ��  5�  �T  5�  �T  5(  ��  5(      H   ,  �<  4`  �<  5(  �  5(  �  4`  �<  4`      H   ,  ��  7�  ��  8H  �t  8H  �t  7�  ��  7�      H   ,  �t  @�  �t  A�  �<  A�  �<  @�  �t  @�      H   ,  �L  5(  �L  5�  �  5�  �  5(  �L  5(      H   ,  �t  7�  �t  8H  �<  8H  �<  7�  �t  7�      H   ,  �4  5�  �4  6�  ��  6�  ��  5�  �4  5�      H   ,  ��  6�  ��  7�  �t  7�  �t  6�  ��  6�      H   ,  �T  4`  �T  5(  �  5(  �  4`  �T  4`      H   ,  ��  5�  ��  6�  ��  6�  ��  5�  ��  5�      H   ,  ��  4`  ��  5(  �T  5(  �T  4`  ��  4`      H   ,  ��  5�  ��  6�  ��  6�  ��  5�  ��  5�      H   ,  ��  5(  ��  5�  ��  5�  ��  5(  ��  5(      H   ,  ��  5�  ��  6�  �t  6�  �t  5�  ��  5�      H   ,  �t  5(  �t  5�  �<  5�  �<  5(  �t  5(      H   ,  ��  5(  ��  5�  ��  5�  ��  5(  ��  5(      H   ,  ��  5(  ��  5�  �t  5�  �t  5(  ��  5(      H   ,  ��  5(  ��  5�  �L  5�  �L  5(  ��  5(      H   ,  ��  5(  ��  5�  ��  5�  ��  5(  ��  5(      H   ,  ��  5(  ��  5�  ��  5�  ��  5(  ��  5(      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  �t  6�  �t  7�  �<  7�  �<  6�  �t  6�      H   ,  �<  8H  �<  9  �  9  �  8H  �<  8H      H   ,  ��  4`  ��  5(  �t  5(  �t  4`  ��  4`      H   ,  �T  6�  �T  7�  �  7�  �  6�  �T  6�      H   ,  ��  6�  ��  7�  ��  7�  ��  6�  ��  6�      H   ,  ��  4`  ��  5(  �L  5(  �L  4`  ��  4`      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  �  7�  �  8H  ��  8H  ��  7�  �  7�      H   ,  �<  5�  �<  6�  �  6�  �  5�  �<  5�      H   ,  �l  4`  �l  5(  �4  5(  �4  4`  �l  4`      H   ,  �t  5�  �t  6�  �<  6�  �<  5�  �t  5�      H   ,  �  6�  �  7�  ��  7�  ��  6�  �  6�      H   ,  ��  5(  ��  5�  ��  5�  ��  5(  ��  5(      H   ,  �<  6�  �<  7�  �  7�  �  6�  �<  6�      H   ,  �  5�  �  6�  ��  6�  ��  5�  �  5�      H   ,  ��  5(  ��  5�  �l  5�  �l  5(  ��  5(      H   ,  �t  4`  �t  5(  �<  5(  �<  4`  �t  4`      H   ,  ��  7�  ��  8H  ��  8H  ��  7�  ��  7�      H   ,  �t  8H  �t  9  �<  9  �<  8H  �t  8H      H   ,  �  5(  �  5�  ��  5�  ��  5(  �  5(      H   ,  �  4`  �  5(  ��  5(  ��  4`  �  4`      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  &P  ��  '  ��  '  ��  &P  ��  &P      H   ,  ��  &P  ��  '  �L  '  �L  &P  ��  &P      H   ,  ��  *8  ��  +   ��  +   ��  *8  ��  *8      H   ,  ��  0x  ��  1@  �L  1@  �L  0x  ��  0x      H   ,  �T  2�  �T  3�  �  3�  �  2�  �T  2�      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  �L  '�  �L  (�  �  (�  �  '�  �L  '�      H   ,  ��  +�  ��  ,�  �L  ,�  �L  +�  ��  +�      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  �L  )p  �L  *8  �  *8  �  )p  �L  )p      H   ,  �l  2  �l  2�  �4  2�  �4  2  �l  2      H   ,  �L  2  �L  2�  �  2�  �  2  �L  2      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  )p  ��  *8  ��  *8  ��  )p  ��  )p      H   ,  ��  +   ��  +�  �L  +�  �L  +   ��  +       H   ,  ��  -X  ��  .   ��  .   ��  -X  ��  -X      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  *8  ��  +   �L  +   �L  *8  ��  *8      H   ,  �L  1@  �L  2  �  2  �  1@  �L  1@      H   ,  ��  ,�  ��  -X  ��  -X  ��  ,�  ��  ,�      H   ,  ��  2  ��  2�  �l  2�  �l  2  ��  2      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  �  2�  �  3�  ��  3�  ��  2�  �  2�      H   ,  ��  )p  ��  *8  �L  *8  �L  )p  ��  )p      H   ,  ��  (�  ��  )p  ��  )p  ��  (�  ��  (�      H   ,  �l  2�  �l  3�  �4  3�  �4  2�  �l  2�      H   ,  �4  2  �4  2�  ��  2�  ��  2  �4  2      H   ,  ��  2�  ��  3�  �L  3�  �L  2�  ��  2�      H   ,  �L  (�  �L  )p  �  )p  �  (�  �L  (�      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  �L  '  �L  '�  �  '�  �  '  �L  '      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  '�  ��  (�  ��  (�  ��  '�  ��  '�      H   ,  �  2�  �  3�  ��  3�  ��  2�  �  2�      H   ,  ��  (�  ��  )p  �L  )p  �L  (�  ��  (�      H   ,  ��  +�  ��  ,�  ��  ,�  ��  +�  ��  +�      H   ,  �  2  �  2�  ��  2�  ��  2  �  2      H   ,  ��  2�  ��  3�  �T  3�  �T  2�  ��  2�      H   ,  ��  2�  ��  3�  �l  3�  �l  2�  ��  2�      H   ,  ��  1@  ��  2  �l  2  �l  1@  ��  1@      H   ,  ��  2  ��  2�  �L  2�  �L  2  ��  2      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  '�  ��  (�  �L  (�  �L  '�  ��  '�      H   ,  �  1@  �  2  ��  2  ��  1@  �  1@      H   ,  ��  2  ��  2�  �T  2�  �T  2  ��  2      H   ,  �L  2�  �L  3�  �  3�  �  2�  �L  2�      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  �L  0x  �L  1@  �  1@  �  0x  �L  0x      H   ,  �L  &P  �L  '  �  '  �  &P  �L  &P      H   ,  �  &P  �  '  ��  '  ��  &P  �  &P      H   ,  ��  '  ��  '�  ��  '�  ��  '  ��  '      H   ,  �4  2�  �4  3�  ��  3�  ��  2�  �4  2�      H   ,  �l  1@  �l  2  �4  2  �4  1@  �l  1@      H   ,  ��  1@  ��  2  �L  2  �L  1@  ��  1@      H   ,  ��  +   ��  +�  ��  +�  ��  +   ��  +       H   ,  ��  '  ��  '�  �L  '�  �L  '  ��  '      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  �|  3�  �|  4`  �D  4`  �D  3�  �|  3�      H   ,  ��  5(  ��  5�  �t  5�  �t  5(  ��  5(      H   ,  ��  8H  ��  9  �t  9  �t  8H  ��  8H      H   ,  ��  4`  ��  5(  �t  5(  �t  4`  ��  4`      H   ,  �T  3�  �T  4`  �  4`  �  3�  �T  3�      H   ,  ��  9  ��  9�  �t  9�  �t  9  ��  9      H   ,  ��  3�  ��  4`  �t  4`  �t  3�  ��  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  ��  2�  ��  3�  �t  3�  �t  2�  ��  2�      H   ,  �$  3�  �$  4`  ��  4`  ��  3�  �$  3�      H   ,  �t  3�  �t  4`  �<  4`  �<  3�  �t  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  ��  2  ��  2�  �t  2�  �t  2  ��  2      H   ,  ��  3�  ��  4`  �|  4`  �|  3�  ��  3�      H   ,  ��  1@  ��  2  �t  2  �t  1@  ��  1@      H   ,  ��  7�  ��  8H  �t  8H  �t  7�  ��  7�      H   ,  �D  3�  �D  4`  �  4`  �  3�  �D  3�      H   ,  ��  0x  ��  1@  �t  1@  �t  0x  ��  0x      H   ,  ��  /�  ��  0x  �t  0x  �t  /�  ��  /�      H   ,  ��  3�  ��  4`  �\  4`  �\  3�  ��  3�      H   ,  ��  6�  ��  7�  �t  7�  �t  6�  ��  6�      H   ,  ��  .�  ��  /�  �t  /�  �t  .�  ��  .�      H   ,  �\  3�  �\  4`  �$  4`  �$  3�  �\  3�      H   ,  ��  3�  ��  4`  �d  4`  �d  3�  ��  3�      H   ,  �  3�  �  4`  ��  4`  ��  3�  �  3�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  �  3�  �  4`  ��  4`  ��  3�  �  3�      H   ,  �,  3�  �,  4`  ��  4`  ��  3�  �,  3�      H   ,  ��  5�  ��  6�  �t  6�  �t  5�  ��  5�      H   ,  ��  3�  ��  4`  ��  4`  ��  3�  ��  3�      H   ,  ��  ;h  ��  <0  �t  <0  �t  ;h  ��  ;h      H   ,  �d  3�  �d  4`  �,  4`  �,  3�  �d  3�      H   ,  ��  :�  ��  ;h  �t  ;h  �t  :�  ��  :�      H   ,  ��  9�  ��  :�  �t  :�  �t  9�  ��  9�      H   ,  ��  3�  ��  4`  �T  4`  �T  3�  ��  3�      H   ,  ��  :�  ��  ;h  ��  ;h  ��  :�  ��  :�      H   ,  ��  4`  ��  5(  �|  5(  �|  4`  ��  4`      H   ,  �$  :�  �$  ;h  ��  ;h  ��  :�  �$  :�      H   ,  ��  8H  ��  9  �|  9  �|  8H  ��  8H      H   ,  ��  :�  ��  ;h  �\  ;h  �\  :�  ��  :�      H   ,  �  :�  �  ;h  ��  ;h  ��  :�  �  :�      H   ,  ��  5�  ��  6�  �|  6�  �|  5�  ��  5�      H   ,  �<  :�  �<  ;h  �  ;h  �  :�  �<  :�      H   ,  �|  :�  �|  ;h  �D  ;h  �D  :�  �|  :�      H   ,  ��  9  ��  9�  �|  9�  �|  9  ��  9      H   ,  ��  7�  ��  8H  �|  8H  �|  7�  ��  7�      H   ,  ��  @�  ��  A�  �|  A�  �|  @�  ��  @�      H   ,  ��  @  ��  @�  �|  @�  �|  @  ��  @      H   ,  �D  :�  �D  ;h  �  ;h  �  :�  �D  :�      H   ,  ��  >�  ��  ?P  �|  ?P  �|  >�  ��  >�      H   ,  ��  =�  ��  >�  �|  >�  �|  =�  ��  =�      H   ,  ��  <�  ��  =�  �|  =�  �|  <�  ��  <�      H   ,  ��  :�  ��  ;h  ��  ;h  ��  :�  ��  :�      H   ,  ��  <0  ��  <�  �|  <�  �|  <0  ��  <0      H   ,  ��  5(  ��  5�  �|  5�  �|  5(  ��  5(      H   ,  ��  ;h  ��  <0  �|  <0  �|  ;h  ��  ;h      H   ,  �t  :�  �t  ;h  �<  ;h  �<  :�  �t  :�      H   ,  ��  6�  ��  7�  �|  7�  �|  6�  ��  6�      H   ,  ��  :�  ��  ;h  �|  ;h  �|  :�  ��  :�      H   ,  �\  :�  �\  ;h  �$  ;h  �$  :�  �\  :�      H   ,  ��  9�  ��  :�  �|  :�  �|  9�  ��  9�      H   ,  �D  ;h  �D  <0  �  <0  �  ;h  �D  ;h      H   ,  �|  <0  �|  <�  �D  <�  �D  <0  �|  <0      H   ,  �|  <�  �|  =�  �D  =�  �D  <�  �|  <�      H   ,  �|  ;h  �|  <0  �D  <0  �D  ;h  �|  ;h      H   ,  ��  >�  ��  ?P  ��  ?P  ��  >�  ��  >�      H   ,  �$  <�  �$  =�  ��  =�  ��  <�  �$  <�      H   ,  �  <0  �  <�  ��  <�  ��  <0  �  <0      H   ,  ��  @�  ��  A�  �\  A�  �\  @�  ��  @�      H   ,  ��  <�  ��  =�  ��  =�  ��  <�  ��  <�      H   ,  ��  =�  ��  >�  ��  >�  ��  =�  ��  =�      H   ,  �<  @  �<  @�  �  @�  �  @  �<  @      H   ,  ��  ?P  ��  @  �\  @  �\  ?P  ��  ?P      H   ,  ��  <�  ��  =�  ��  =�  ��  <�  ��  <�      H   ,  ��  <�  ��  =�  �\  =�  �\  <�  ��  <�      H   ,  �  ;h  �  <0  ��  <0  ��  ;h  �  ;h      H   ,  ��  =�  ��  >�  ��  >�  ��  =�  ��  =�      H   ,  �  @�  �  A�  ��  A�  ��  @�  �  @�      H   ,  �$  <0  �$  <�  ��  <�  ��  <0  �$  <0      H   ,  �$  >�  �$  ?P  ��  ?P  ��  >�  �$  >�      H   ,  ��  @�  ��  A�  ��  A�  ��  @�  ��  @�      H   ,  ��  ;h  ��  <0  ��  <0  ��  ;h  ��  ;h      H   ,  ��  <0  ��  <�  �\  <�  �\  <0  ��  <0      H   ,  �$  @  �$  @�  ��  @�  ��  @  �$  @      H   ,  ��  <0  ��  <�  ��  <�  ��  <0  ��  <0      H   ,  �<  ;h  �<  <0  �  <0  �  ;h  �<  ;h      H   ,  �<  <�  �<  =�  �  =�  �  <�  �<  <�      H   ,  �\  @�  �\  A�  �$  A�  �$  @�  �\  @�      H   ,  ��  @  ��  @�  ��  @�  ��  @  ��  @      H   ,  �\  @  �\  @�  �$  @�  �$  @  �\  @      H   ,  �  <�  �  =�  ��  =�  ��  <�  �  <�      H   ,  �<  =�  �<  >�  �  >�  �  =�  �<  =�      H   ,  �  @  �  @�  ��  @�  ��  @  �  @      H   ,  �t  <�  �t  =�  �<  =�  �<  <�  �t  <�      H   ,  �\  ?P  �\  @  �$  @  �$  ?P  �\  ?P      H   ,  ��  =�  ��  >�  �\  >�  �\  =�  ��  =�      H   ,  ��  ;h  ��  <0  �\  <0  �\  ;h  ��  ;h      H   ,  �t  <0  �t  <�  �<  <�  �<  <0  �t  <0      H   ,  �\  >�  �\  ?P  �$  ?P  �$  >�  �\  >�      H   ,  �<  >�  �<  ?P  �  ?P  �  >�  �<  >�      H   ,  ��  >�  ��  ?P  �\  ?P  �\  >�  ��  >�      H   ,  ��  ?P  ��  @  ��  @  ��  ?P  ��  ?P      H   ,  �$  ;h  �$  <0  ��  <0  ��  ;h  �$  ;h      H   ,  �t  ;h  �t  <0  �<  <0  �<  ;h  �t  ;h      H   ,  �\  =�  �\  >�  �$  >�  �$  =�  �\  =�      H   ,  ��  <0  ��  <�  ��  <�  ��  <0  ��  <0      H   ,  �  =�  �  >�  ��  >�  ��  =�  �  =�      H   ,  ��  @�  ��  A�  ��  A�  ��  @�  ��  @�      H   ,  �$  =�  �$  >�  ��  >�  ��  =�  �$  =�      H   ,  �  >�  �  ?P  ��  ?P  ��  >�  �  >�      H   ,  �\  <�  �\  =�  �$  =�  �$  <�  �\  <�      H   ,  �<  <0  �<  <�  �  <�  �  <0  �<  <0      H   ,  �  ?P  �  @  ��  @  ��  ?P  �  ?P      H   ,  �\  <0  �\  <�  �$  <�  �$  <0  �\  <0      H   ,  ��  >�  ��  ?P  ��  ?P  ��  >�  ��  >�      H   ,  ��  @  ��  @�  ��  @�  ��  @  ��  @      H   ,  �$  @�  �$  A�  ��  A�  ��  @�  �$  @�      H   ,  �\  ;h  �\  <0  �$  <0  �$  ;h  �\  ;h      H   ,  �<  @�  �<  A�  �  A�  �  @�  �<  @�      H   ,  ��  @  ��  @�  �\  @�  �\  @  ��  @      H   ,  ��  ?P  ��  @  ��  @  ��  ?P  ��  ?P      H   ,  ��  ;h  ��  <0  ��  <0  ��  ;h  ��  ;h      H   ,  �$  ?P  �$  @  ��  @  ��  ?P  �$  ?P      H   ,  ��  8H  ��  9  ��  9  ��  8H  ��  8H      H   ,  ��  6�  ��  7�  ��  7�  ��  6�  ��  6�      H   ,  ��  8H  ��  9  ��  9  ��  8H  ��  8H      H   ,  �t  5�  �t  6�  �<  6�  �<  5�  �t  5�      H   ,  �  9�  �  :�  ��  :�  ��  9�  �  9�      H   ,  ��  9�  ��  :�  ��  :�  ��  9�  ��  9�      H   ,  �  7�  �  8H  ��  8H  ��  7�  �  7�      H   ,  ��  9  ��  9�  ��  9�  ��  9  ��  9      H   ,  �t  5(  �t  5�  �<  5�  �<  5(  �t  5(      H   ,  ��  9  ��  9�  �\  9�  �\  9  ��  9      H   ,  �<  9�  �<  :�  �  :�  �  9�  �<  9�      H   ,  �$  9  �$  9�  ��  9�  ��  9  �$  9      H   ,  �$  9�  �$  :�  ��  :�  ��  9�  �$  9�      H   ,  �<  7�  �<  8H  �  8H  �  7�  �<  7�      H   ,  �\  9  �\  9�  �$  9�  �$  9  �\  9      H   ,  �<  5(  �<  5�  �  5�  �  5(  �<  5(      H   ,  �<  5�  �<  6�  �  6�  �  5�  �<  5�      H   ,  �  6�  �  7�  ��  7�  ��  6�  �  6�      H   ,  �  9  �  9�  ��  9�  ��  9  �  9      H   ,  �<  8H  �<  9  �  9  �  8H  �<  8H      H   ,  ��  5�  ��  6�  ��  6�  ��  5�  ��  5�      H   ,  ��  7�  ��  8H  ��  8H  ��  7�  ��  7�      H   ,  �t  9�  �t  :�  �<  :�  �<  9�  �t  9�      H   ,  �<  4`  �<  5(  �  5(  �  4`  �<  4`      H   ,  ��  9�  ��  :�  ��  :�  ��  9�  ��  9�      H   ,  �  5�  �  6�  ��  6�  ��  5�  �  5�      H   ,  �$  7�  �$  8H  ��  8H  ��  7�  �$  7�      H   ,  �t  9  �t  9�  �<  9�  �<  9  �t  9      H   ,  ��  9  ��  9�  ��  9�  ��  9  ��  9      H   ,  �<  6�  �<  7�  �  7�  �  6�  �<  6�      H   ,  ��  9�  ��  :�  �\  :�  �\  9�  ��  9�      H   ,  �t  6�  �t  7�  �<  7�  �<  6�  �t  6�      H   ,  �t  8H  �t  9  �<  9  �<  8H  �t  8H      H   ,  �<  9  �<  9�  �  9�  �  9  �<  9      H   ,  �$  8H  �$  9  ��  9  ��  8H  �$  8H      H   ,  �t  4`  �t  5(  �<  5(  �<  4`  �t  4`      H   ,  �  8H  �  9  ��  9  ��  8H  �  8H      H   ,  ��  7�  ��  8H  ��  8H  ��  7�  ��  7�      H   ,  �t  7�  �t  8H  �<  8H  �<  7�  �t  7�      H   ,  �\  9�  �\  :�  �$  :�  �$  9�  �\  9�      H   ,  �|  7�  �|  8H  �D  8H  �D  7�  �|  7�      H   ,  �D  7�  �D  8H  �  8H  �  7�  �D  7�      H   ,  �D  6�  �D  7�  �  7�  �  6�  �D  6�      H   ,  �D  9�  �D  :�  �  :�  �  9�  �D  9�      H   ,  ��  5�  ��  6�  �d  6�  �d  5�  ��  5�      H   ,  �  5�  �  6�  ��  6�  ��  5�  �  5�      H   ,  �d  4`  �d  5(  �,  5(  �,  4`  �d  4`      H   ,  �|  9�  �|  :�  �D  :�  �D  9�  �|  9�      H   ,  �D  8H  �D  9  �  9  �  8H  �D  8H      H   ,  �  4`  �  5(  ��  5(  ��  4`  �  4`      H   ,  ��  8H  ��  9  ��  9  ��  8H  ��  8H      H   ,  �  5(  �  5�  ��  5�  ��  5(  �  5(      H   ,  ��  5(  ��  5�  �d  5�  �d  5(  ��  5(      H   ,  �D  9  �D  9�  �  9�  �  9  �D  9      H   ,  �|  8H  �|  9  �D  9  �D  8H  �|  8H      H   ,  �|  6�  �|  7�  �D  7�  �D  6�  �|  6�      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  �D  5�  �D  6�  �  6�  �  5�  �D  5�      H   ,  �,  4`  �,  5(  ��  5(  ��  4`  �,  4`      H   ,  �D  4`  �D  5(  �  5(  �  4`  �D  4`      H   ,  �  7�  �  8H  ��  8H  ��  7�  �  7�      H   ,  �|  5(  �|  5�  �D  5�  �D  5(  �|  5(      H   ,  �  8H  �  9  ��  9  ��  8H  �  8H      H   ,  ��  4`  ��  5(  �d  5(  �d  4`  ��  4`      H   ,  �  9�  �  :�  ��  :�  ��  9�  �  9�      H   ,  �|  4`  �|  5(  �D  5(  �D  4`  �|  4`      H   ,  ��  5(  ��  5�  ��  5�  ��  5(  ��  5(      H   ,  ��  7�  ��  8H  ��  8H  ��  7�  ��  7�      H   ,  ��  6�  ��  7�  ��  7�  ��  6�  ��  6�      H   ,  �D  5(  �D  5�  �  5�  �  5(  �D  5(      H   ,  �|  9  �|  9�  �D  9�  �D  9  �|  9      H   ,  ��  5�  ��  6�  ��  6�  ��  5�  ��  5�      H   ,  �|  5�  �|  6�  �D  6�  �D  5�  �|  5�      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  �  6�  �  7�  ��  7�  ��  6�  �  6�      H   ,  �  9  �  9�  ��  9�  ��  9  �  9      H   ,  ��  8H  ��  9  ��  9  ��  8H  ��  8H      H   ,  �T  4`  �T  5(  �  5(  �  4`  �T  4`      H   ,  �  7�  �  8H  ��  8H  ��  7�  �  7�      H   ,  ��  5�  ��  6�  ��  6�  ��  5�  ��  5�      H   ,  ��  5(  ��  5�  �T  5�  �T  5(  ��  5(      H   ,  �  8H  �  9  ��  9  ��  8H  �  8H      H   ,  �T  5�  �T  6�  �  6�  �  5�  �T  5�      H   ,  ��  9  ��  9�  ��  9�  ��  9  ��  9      H   ,  �T  6�  �T  7�  �  7�  �  6�  �T  6�      H   ,  ��  9�  ��  :�  ��  :�  ��  9�  ��  9�      H   ,  ��  4`  ��  5(  �T  5(  �T  4`  ��  4`      H   ,  ��  6�  ��  7�  ��  7�  ��  6�  ��  6�      H   ,  ��  4`  ��  5(  ��  5(  ��  4`  ��  4`      H   ,  �  5�  �  6�  ��  6�  ��  5�  �  5�      H   ,  ��  7�  ��  8H  ��  8H  ��  7�  ��  7�      H   ,  �  4`  �  5(  ��  5(  ��  4`  �  4`      H   ,  �  5(  �  5�  ��  5�  ��  5(  �  5(      H   ,  ��  5(  ��  5�  ��  5�  ��  5(  ��  5(      H   ,  �T  5(  �T  5�  �  5�  �  5(  �T  5(      H   ,  �  6�  �  7�  ��  7�  ��  6�  �  6�      H   ,  ��  &P  ��  '  �l  '  �l  &P  ��  &P      H   ,  ��  ,�  ��  -X  ��  -X  ��  ,�  ��  ,�      H   ,  ��  *8  ��  +   �l  +   �l  *8  ��  *8      H   ,  ��  )p  ��  *8  �l  *8  �l  )p  ��  )p      H   ,  ��  2  ��  2�  �l  2�  �l  2  ��  2      H   ,  ��  .   ��  .�  �l  .�  �l  .   ��  .       H   ,  ��  -X  ��  .   �l  .   �l  -X  ��  -X      H   ,  ��  .�  ��  /�  �l  /�  �l  .�  ��  .�      H   ,  �l  ,�  �l  -X  �4  -X  �4  ,�  �l  ,�      H   ,  ��  1@  ��  2  �l  2  �l  1@  ��  1@      H   ,  ��  ,�  ��  -X  �l  -X  �l  ,�  ��  ,�      H   ,  ��  ,�  ��  -X  �T  -X  �T  ,�  ��  ,�      H   ,  ��  ,�  ��  -X  ��  -X  ��  ,�  ��  ,�      H   ,  ��  '  ��  '�  �l  '�  �l  '  ��  '      H   ,  ��  +   ��  +�  �l  +�  �l  +   ��  +       H   ,  ��  (�  ��  )p  �l  )p  �l  (�  ��  (�      H   ,  ��  ,�  ��  -X  ��  -X  ��  ,�  ��  ,�      H   ,  ��  /�  ��  0x  �l  0x  �l  /�  ��  /�      H   ,  ��  '�  ��  (�  �l  (�  �l  '�  ��  '�      H   ,  �4  ,�  �4  -X  ��  -X  ��  ,�  �4  ,�      H   ,  ��  +�  ��  ,�  �l  ,�  �l  +�  ��  +�      H   ,  ��  0x  ��  1@  �l  1@  �l  0x  ��  0x      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  .   ��  .�  �T  .�  �T  .   ��  .       H   ,  �  .�  �  /�  ��  /�  ��  .�  �  .�      H   ,  �l  0x  �l  1@  �4  1@  �4  0x  �l  0x      H   ,  �T  -X  �T  .   �  .   �  -X  �T  -X      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �T  /�  �T  0x  �  0x  �  /�  �T  /�      H   ,  �4  1@  �4  2  ��  2  ��  1@  �4  1@      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �l  1@  �l  2  �4  2  �4  1@  �l  1@      H   ,  �T  .�  �T  /�  �  /�  �  .�  �T  .�      H   ,  �4  -X  �4  .   ��  .   ��  -X  �4  -X      H   ,  �  1@  �  2  ��  2  ��  1@  �  1@      H   ,  �  0x  �  1@  ��  1@  ��  0x  �  0x      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  ��  1@  ��  2  �T  2  �T  1@  ��  1@      H   ,  �4  0x  �4  1@  ��  1@  ��  0x  �4  0x      H   ,  ��  2  ��  2�  �T  2�  �T  2  ��  2      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  �T  1@  �T  2  �  2  �  1@  �T  1@      H   ,  �l  /�  �l  0x  �4  0x  �4  /�  �l  /�      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  -X  ��  .   ��  .   ��  -X  ��  -X      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  �4  /�  �4  0x  ��  0x  ��  /�  �4  /�      H   ,  �  2  �  2�  ��  2�  ��  2  �  2      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  ��  2�  ��  3�  �T  3�  �T  2�  ��  2�      H   ,  �l  -X  �l  .   �4  .   �4  -X  �l  -X      H   ,  �T  2�  �T  3�  �  3�  �  2�  �T  2�      H   ,  ��  .�  ��  /�  �T  /�  �T  .�  ��  .�      H   ,  �T  .   �T  .�  �  .�  �  .   �T  .       H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  �l  .�  �l  /�  �4  /�  �4  .�  �l  .�      H   ,  �4  .�  �4  /�  ��  /�  ��  .�  �4  .�      H   ,  �T  0x  �T  1@  �  1@  �  0x  �T  0x      H   ,  �  /�  �  0x  ��  0x  ��  /�  �  /�      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  ��  -X  ��  .   ��  .   ��  -X  ��  -X      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  -X  ��  .   �T  .   �T  -X  ��  -X      H   ,  �4  2  �4  2�  ��  2�  ��  2  �4  2      H   ,  ��  /�  ��  0x  �T  0x  �T  /�  ��  /�      H   ,  �l  2  �l  2�  �4  2�  �4  2  �l  2      H   ,  �  2�  �  3�  ��  3�  ��  2�  �  2�      H   ,  ��  0x  ��  1@  �T  1@  �T  0x  ��  0x      H   ,  �4  .   �4  .�  ��  .�  ��  .   �4  .       H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  �T  2  �T  2�  �  2�  �  2  �T  2      H   ,  �l  .   �l  .�  �4  .�  �4  .   �l  .       H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  �L  0x  �L  1@  �  1@  �  0x  �L  0x      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  0x  ��  1@  �L  1@  �L  0x  ��  0x      H   ,  �,  1@  �,  2  ��  2  ��  1@  �,  1@      H   ,  �  /�  �  0x  ��  0x  ��  /�  �  /�      H   ,  �L  .   �L  .�  �  .�  �  .   �L  .       H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �,  .�  �,  /�  ��  /�  ��  .�  �,  .�      H   ,  �d  /�  �d  0x  �,  0x  �,  /�  �d  /�      H   ,  �d  1@  �d  2  �,  2  �,  1@  �d  1@      H   ,  �  1@  �  2  ��  2  ��  1@  �  1@      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �,  0x  �,  1@  ��  1@  ��  0x  �,  0x      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  2  ��  2�  �L  2�  �L  2  ��  2      H   ,  �L  .�  �L  /�  �  /�  �  .�  �L  .�      H   ,  �,  .   �,  .�  ��  .�  ��  .   �,  .       H   ,  ��  .   ��  .�  �L  .�  �L  .   ��  .       H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �  2  �  2�  ��  2�  ��  2  �  2      H   ,  �d  .�  �d  /�  �,  /�  �,  .�  �d  .�      H   ,  �  .�  �  /�  ��  /�  ��  .�  �  .�      H   ,  �,  2  �,  2�  ��  2�  ��  2  �,  2      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �  .   �  .�  ��  .�  ��  .   �  .       H   ,  �L  2  �L  2�  �  2�  �  2  �L  2      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  ��  /�  ��  0x  �L  0x  �L  /�  ��  /�      H   ,  �d  2  �d  2�  �,  2�  �,  2  �d  2      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  �d  .   �d  .�  �,  .�  �,  .   �d  .       H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  .�  ��  /�  �L  /�  �L  .�  ��  .�      H   ,  �,  /�  �,  0x  ��  0x  ��  /�  �,  /�      H   ,  �d  0x  �d  1@  �,  1@  �,  0x  �d  0x      H   ,  �  0x  �  1@  ��  1@  ��  0x  �  0x      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  1@  ��  2  �L  2  �L  1@  ��  1@      H   ,  �L  1@  �L  2  �  2  �  1@  �L  1@      H   ,  �L  /�  �L  0x  �  0x  �  /�  �L  /�      H   ,  ��  &P  ��  '  ��  '  ��  &P  ��  &P      H   ,  �  *8  �  +   ��  +   ��  *8  �  *8      H   ,  ��  '  ��  '�  �L  '�  �L  '  ��  '      H   ,  ��  (�  ��  )p  ��  )p  ��  (�  ��  (�      H   ,  ��  *8  ��  +   ��  +   ��  *8  ��  *8      H   ,  ��  &P  ��  '  ��  '  ��  &P  ��  &P      H   ,  �  +�  �  ,�  ��  ,�  ��  +�  �  +�      H   ,  ��  (�  ��  )p  �L  )p  �L  (�  ��  (�      H   ,  �L  )p  �L  *8  �  *8  �  )p  �L  )p      H   ,  �  +   �  +�  ��  +�  ��  +   �  +       H   ,  �  (�  �  )p  ��  )p  ��  (�  �  (�      H   ,  �L  &P  �L  '  �  '  �  &P  �L  &P      H   ,  ��  &P  ��  '  �L  '  �L  &P  ��  &P      H   ,  ��  +�  ��  ,�  ��  ,�  ��  +�  ��  +�      H   ,  �  &P  �  '  ��  '  ��  &P  �  &P      H   ,  ��  '  ��  '�  ��  '�  ��  '  ��  '      H   ,  �L  *8  �L  +   �  +   �  *8  �L  *8      H   ,  �d  &P  �d  '  �,  '  �,  &P  �d  &P      H   ,  ��  '�  ��  (�  �L  (�  �L  '�  ��  '�      H   ,  ��  )p  ��  *8  ��  *8  ��  )p  ��  )p      H   ,  ��  '�  ��  (�  ��  (�  ��  '�  ��  '�      H   ,  �  )p  �  *8  ��  *8  ��  )p  �  )p      H   ,  ��  '  ��  '�  ��  '�  ��  '  ��  '      H   ,  ��  '�  ��  (�  ��  (�  ��  '�  ��  '�      H   ,  ��  +   ��  +�  ��  +�  ��  +   ��  +       H   ,  �  '  �  '�  ��  '�  ��  '  �  '      H   ,  �  '�  �  (�  ��  (�  ��  '�  �  '�      H   ,  ��  &P  ��  '  ��  '  ��  &P  ��  &P      H   ,  �L  '  �L  '�  �  '�  �  '  �L  '      H   ,  �L  '�  �L  (�  �  (�  �  '�  �L  '�      H   ,  �L  (�  �L  )p  �  )p  �  (�  �L  (�      H   ,  �l  '  �l  '�  �4  '�  �4  '  �l  '      H   ,  �l  &P  �l  '  �4  '  �4  &P  �l  &P      H   ,  ��  *8  ��  +   ��  +   ��  *8  ��  *8      H   ,  �4  +   �4  +�  ��  +�  ��  +   �4  +       H   ,  �4  )p  �4  *8  ��  *8  ��  )p  �4  )p      H   ,  ��  +�  ��  ,�  �T  ,�  �T  +�  ��  +�      H   ,  �4  *8  �4  +   ��  +   ��  *8  �4  *8      H   ,  �4  +�  �4  ,�  ��  ,�  ��  +�  �4  +�      H   ,  ��  +   ��  +�  ��  +�  ��  +   ��  +       H   ,  �l  +   �l  +�  �4  +�  �4  +   �l  +       H   ,  ��  +�  ��  ,�  ��  ,�  ��  +�  ��  +�      H   ,  �l  +�  �l  ,�  �4  ,�  �4  +�  �l  +�      H   ,  �l  (�  �l  )p  �4  )p  �4  (�  �l  (�      H   ,  �l  '�  �l  (�  �4  (�  �4  '�  �l  '�      H   ,  ��  )p  ��  *8  ��  *8  ��  )p  ��  )p      H   ,  �l  )p  �l  *8  �4  *8  �4  )p  �l  )p      H   ,  ��  +�  ��  ,�  ��  ,�  ��  +�  ��  +�      H   ,  ��  +   ��  +�  ��  +�  ��  +   ��  +       H   ,  �4  (�  �4  )p  ��  )p  ��  (�  �4  (�      H   ,  �4  '�  �4  (�  ��  (�  ��  '�  �4  '�      H   ,  �l  *8  �l  +   �4  +   �4  *8  �l  *8      H   ,  ��  *8  ��  +   ��  +   ��  *8  ��  *8      H   ,  �d  ,�  �d  -X  �,  -X  �,  ,�  �d  ,�      H   ,  ��  ,�  ��  -X  ��  -X  ��  ,�  ��  ,�      H   ,  ��  ,�  ��  -X  �d  -X  �d  ,�  ��  ,�      H   ,  ��  /�  ��  0x  �|  0x  �|  /�  ��  /�      H   ,  ��  2�  ��  3�  �|  3�  �|  2�  ��  2�      H   ,  ��  1@  ��  2  �|  2  �|  1@  ��  1@      H   ,  ��  ,�  ��  -X  ��  -X  ��  ,�  ��  ,�      H   ,  ��  0x  ��  1@  �|  1@  �|  0x  ��  0x      H   ,  �,  ,�  �,  -X  ��  -X  ��  ,�  �,  ,�      H   ,  ��  2  ��  2�  �|  2�  �|  2  ��  2      H   ,  ��  2  ��  2�  �d  2�  �d  2  ��  2      H   ,  �  /�  �  0x  ��  0x  ��  /�  �  /�      H   ,  �d  -X  �d  .   �,  .   �,  -X  �d  -X      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �  1@  �  2  ��  2  ��  1@  �  1@      H   ,  �|  2  �|  2�  �D  2�  �D  2  �|  2      H   ,  �|  1@  �|  2  �D  2  �D  1@  �|  1@      H   ,  �D  0x  �D  1@  �  1@  �  0x  �D  0x      H   ,  �D  1@  �D  2  �  2  �  1@  �D  1@      H   ,  �d  .�  �d  /�  �,  /�  �,  .�  �d  .�      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  ��  1@  ��  2  �d  2  �d  1@  ��  1@      H   ,  �,  2�  �,  3�  ��  3�  ��  2�  �,  2�      H   ,  �d  /�  �d  0x  �,  0x  �,  /�  �d  /�      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  �d  .   �d  .�  �,  .�  �,  .   �d  .       H   ,  �,  2  �,  2�  ��  2�  ��  2  �,  2      H   ,  �,  -X  �,  .   ��  .   ��  -X  �,  -X      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  �D  2  �D  2�  �  2�  �  2  �D  2      H   ,  �|  0x  �|  1@  �D  1@  �D  0x  �|  0x      H   ,  ��  0x  ��  1@  �d  1@  �d  0x  ��  0x      H   ,  �d  0x  �d  1@  �,  1@  �,  0x  �d  0x      H   ,  �,  1@  �,  2  ��  2  ��  1@  �,  1@      H   ,  �  .�  �  /�  ��  /�  ��  .�  �  .�      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  �  2�  �  3�  ��  3�  ��  2�  �  2�      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  �d  1@  �d  2  �,  2  �,  1@  �d  1@      H   ,  ��  .   ��  .�  �d  .�  �d  .   ��  .       H   ,  �  0x  �  1@  ��  1@  ��  0x  �  0x      H   ,  �,  0x  �,  1@  ��  1@  ��  0x  �,  0x      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  ��  .   ��  .�  ��  .�  ��  .   ��  .       H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  /�  ��  0x  �d  0x  �d  /�  ��  /�      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �|  2�  �|  3�  �D  3�  �D  2�  �|  2�      H   ,  ��  -X  ��  .   �d  .   �d  -X  ��  -X      H   ,  �,  /�  �,  0x  ��  0x  ��  /�  �,  /�      H   ,  �  -X  �  .   ��  .   ��  -X  �  -X      H   ,  �d  2�  �d  3�  �,  3�  �,  2�  �d  2�      H   ,  �D  2�  �D  3�  �  3�  �  2�  �D  2�      H   ,  �  .   �  .�  ��  .�  ��  .   �  .       H   ,  �,  .�  �,  /�  ��  /�  ��  .�  �,  .�      H   ,  �D  /�  �D  0x  �  0x  �  /�  �D  /�      H   ,  �|  /�  �|  0x  �D  0x  �D  /�  �|  /�      H   ,  ��  -X  ��  .   ��  .   ��  -X  ��  -X      H   ,  ��  .�  ��  /�  �d  /�  �d  .�  ��  .�      H   ,  �  2  �  2�  ��  2�  ��  2  �  2      H   ,  �d  2  �d  2�  �,  2�  �,  2  �d  2      H   ,  ��  -X  ��  .   ��  .   ��  -X  ��  -X      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  �,  .   �,  .�  ��  .�  ��  .   �,  .       H   ,  ��  2�  ��  3�  �d  3�  �d  2�  ��  2�      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  �t  2  �t  2�  �<  2�  �<  2  �t  2      H   ,  �$  1@  �$  2  ��  2  ��  1@  �$  1@      H   ,  �<  /�  �<  0x  �  0x  �  /�  �<  /�      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �  .�  �  /�  ��  /�  ��  .�  �  .�      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  ��  .�  ��  /�  ��  /�  ��  .�  ��  .�      H   ,  �$  2�  �$  3�  ��  3�  ��  2�  �$  2�      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  ��  2  ��  2�  �\  2�  �\  2  ��  2      H   ,  �  /�  �  0x  ��  0x  ��  /�  �  /�      H   ,  �t  0x  �t  1@  �<  1@  �<  0x  �t  0x      H   ,  ��  2�  ��  3�  �\  3�  �\  2�  ��  2�      H   ,  �\  .�  �\  /�  �$  /�  �$  .�  �\  .�      H   ,  �<  2  �<  2�  �  2�  �  2  �<  2      H   ,  ��  /�  ��  0x  �\  0x  �\  /�  ��  /�      H   ,  �  2  �  2�  ��  2�  ��  2  �  2      H   ,  �$  2  �$  2�  ��  2�  ��  2  �$  2      H   ,  �\  /�  �\  0x  �$  0x  �$  /�  �\  /�      H   ,  �<  .�  �<  /�  �  /�  �  .�  �<  .�      H   ,  ��  1@  ��  2  ��  2  ��  1@  ��  1@      H   ,  ��  0x  ��  1@  ��  1@  ��  0x  ��  0x      H   ,  �t  1@  �t  2  �<  2  �<  1@  �t  1@      H   ,  ��  2�  ��  3�  ��  3�  ��  2�  ��  2�      H   ,  �  0x  �  1@  ��  1@  ��  0x  �  0x      H   ,  �  1@  �  2  ��  2  ��  1@  �  1@      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  �t  /�  �t  0x  �<  0x  �<  /�  �t  /�      H   ,  �\  2  �\  2�  �$  2�  �$  2  �\  2      H   ,  �\  0x  �\  1@  �$  1@  �$  0x  �\  0x      H   ,  ��  2  ��  2�  ��  2�  ��  2  ��  2      H   ,  �<  2�  �<  3�  �  3�  �  2�  �<  2�      H   ,  �  2�  �  3�  ��  3�  ��  2�  �  2�      H   ,  �$  0x  �$  1@  ��  1@  ��  0x  �$  0x      H   ,  �<  1@  �<  2  �  2  �  1@  �<  1@      H   ,  ��  /�  ��  0x  ��  0x  ��  /�  ��  /�      H   ,  �t  2�  �t  3�  �<  3�  �<  2�  �t  2�      H   ,  ��  .�  ��  /�  �\  /�  �\  .�  ��  .�      H   ,  �t  .�  �t  /�  �<  /�  �<  .�  �t  .�      H   ,  ��  0x  ��  1@  �\  1@  �\  0x  ��  0x      H   ,  ��  1@  ��  2  �\  2  �\  1@  ��  1@      H   ,  �\  1@  �\  2  �$  2  �$  1@  �\  1@      H   ,  �$  .�  �$  /�  ��  /�  ��  .�  �$  .�      H   ,  �$  /�  �$  0x  ��  0x  ��  /�  �$  /�      H   ,  �\  2�  �\  3�  �$  3�  �$  2�  �\  2�      H   ,  �<  0x  �<  1@  �  1@  �  0x  �<  0x      H   ,  ��  *8  ��  +   ��  +   ��  *8  ��  *8      H   ,  ��  +   ��  +�  �d  +�  �d  +   ��  +       H   ,  ��  +�  ��  ,�  ��  ,�  ��  +�  ��  +�      H   ,  �d  +   �d  +�  �,  +�  �,  +   �d  +       H   ,  ��  '  ��  '�  ��  '�  ��  '  ��  '      H   ,  ��  '�  ��  (�  ��  (�  ��  '�  ��  '�      H   ,  �d  (�  �d  )p  �,  )p  �,  (�  �d  (�      H   ,  �,  (�  �,  )p  ��  )p  ��  (�  �,  (�      H   ,  �d  *8  �d  +   �,  +   �,  *8  �d  *8      H   ,  �d  '  �d  '�  �,  '�  �,  '  �d  '      H   ,  ��  +   ��  +�  ��  +�  ��  +   ��  +       H   ,  ��  &P  ��  '  ��  '  ��  &P  ��  &P      H   ,  �,  +   �,  +�  ��  +�  ��  +   �,  +       H   ,  ��  )p  ��  *8  ��  *8  ��  )p  ��  )p      H   ,  �,  )p  �,  *8  ��  *8  ��  )p  �,  )p      H   ,  ��  *8  ��  +   �d  +   �d  *8  ��  *8      H   ,  ��  +�  ��  ,�  ��  ,�  ��  +�  ��  +�      H   ,  �d  +�  �d  ,�  �,  ,�  �,  +�  �d  +�      H   ,  �,  '  �,  '�  ��  '�  ��  '  �,  '      H   ,  �d  '�  �d  (�  �,  (�  �,  '�  �d  '�      H   ,  ��  +�  ��  ,�  �d  ,�  �d  +�  ��  +�      H   ,  �,  '�  �,  (�  ��  (�  ��  '�  �,  '�      H   ,  �d  &P  �d  '  �,  '  �,  &P  �d  &P      H   ,  ��  )p  ��  *8  �d  *8  �d  )p  ��  )p      H   ,  �,  +�  �,  ,�  ��  ,�  ��  +�  �,  +�      H   ,  �,  *8  �,  +   ��  +   ��  *8  �,  *8      H   ,  ��  (�  ��  )p  ��  )p  ��  (�  ��  (�      H   ,  �,  &P  �,  '  ��  '  ��  &P  �,  &P      H   ,  �d  )p  �d  *8  �,  *8  �,  )p  �d  )p      H   ,  ��  8  ��     �t     �t  8  ��  8      H   ,  �T  @  �T    �    �  @  �T  @      H   ,  ��     ��  �  �t  �  �t     ��         H   ,  �  @  �    ��    ��  @  �  @      H   ,  ��  X  ��     �t     �t  X  ��  X      H   ,  �l  @  �l    �4    �4  @  �l  @      H   ,  ��  @  ��    ��    ��  @  ��  @      H   ,  ��  �  ��  X  �t  X  �t  �  ��  �      H   ,  ��  @  ��    ��    ��  @  ��  @      H   ,  ��  �  ��  x  �t  x  �t  �  ��  �      H   ,  ��  @  ��    �l    �l  @  ��  @      H   ,  ��  @  ��    �T    �T  @  ��  @      H   ,  ��  �  ��  �  �t  �  �t  �  ��  �      H   ,  ��  @  ��    ��    ��  @  ��  @      H   ,  ��     ��  �  �t  �  �t     ��         H   ,  ��  �  ��  �  �t  �  �t  �  ��  �      H   ,  �4  @  �4    ��    ��  @  �4  @      H   ,  ��     ��   �  ��   �  ��     ��         H   ,  �,  $�  �,  %�  ��  %�  ��  $�  �,  $�      H   ,  ��   �  ��  !�  ��  !�  ��   �  ��   �      H   ,  ��  $�  ��  %�  ��  %�  ��  $�  ��  $�      H   ,  ��  "h  ��  #0  ��  #0  ��  "h  ��  "h      H   ,  �,  %�  �,  &P  ��  &P  ��  %�  �,  %�      H   ,  �,  #�  �,  $�  ��  $�  ��  #�  �,  #�      H   ,  ��  #0  ��  #�  ��  #�  ��  #0  ��  #0      H   ,  ��  %�  ��  &P  ��  &P  ��  %�  ��  %�      H   ,  ��  #�  ��  $�  ��  $�  ��  #�  ��  #�      H   ,  ��  !�  ��  "h  ��  "h  ��  !�  ��  !�      H   ,  ��  H  ��     �L     �L  H  ��  H      H   ,  ��  H  ��     ��     ��  H  ��  H      H   ,  ��  `  ��  (  �l  (  �l  `  ��  `      H   ,  ��  H  ��     ��     ��  H  ��  H      H   ,  ��  (  ��  �  �l  �  �l  (  ��  (      H   ,  ��  �  ��  `  �l  `  �l  �  ��  �      H   ,  ��  H  ��     ��     ��  H  ��  H      H   ,  ��  %�  ��  &P  �l  &P  �l  %�  ��  %�      H   ,  �,  H  �,     ��     ��  H  �,  H      H   ,  �  H  �     ��     ��  H  �  H      H   ,  ��  �  ��  �  �l  �  �l  �  ��  �      H   ,  ��  �  ��  �  �l  �  �l  �  ��  �      H   ,  �L  H  �L     �     �  H  �L  H      H   ,  ��  �  ��  �  �l  �  �l  �  ��  �      H   ,  �d  H  �d     �,     �,  H  �d  H      H   ,  ��    ��  �  �l  �  �l    ��        H   ,  ��  �  ��  H  �l  H  �l  �  ��  �      H   ,  �d   �  �d  !�  �,  !�  �,   �  �d   �      H   ,  �L  "h  �L  #0  �  #0  �  "h  �L  "h      H   ,  ��   �  ��  !�  ��  !�  ��   �  ��   �      H   ,  �,  #�  �,  $�  ��  $�  ��  #�  �,  #�      H   ,  �  #0  �  #�  ��  #�  ��  #0  �  #0      H   ,  ��  #�  ��  $�  ��  $�  ��  #�  ��  #�      H   ,  �L  #0  �L  #�  �  #�  �  #0  �L  #0      H   ,  �,  !�  �,  "h  ��  "h  ��  !�  �,  !�      H   ,  �,     �,   �  ��   �  ��     �,         H   ,  ��     ��   �  ��   �  ��     ��         H   ,  �,  "h  �,  #0  ��  #0  ��  "h  �,  "h      H   ,  ��  #0  ��  #�  �L  #�  �L  #0  ��  #0      H   ,  �d  !�  �d  "h  �,  "h  �,  !�  �d  !�      H   ,  �     �   �  ��   �  ��     �         H   ,  �d  #0  �d  #�  �,  #�  �,  #0  �d  #0      H   ,  �L  !�  �L  "h  �  "h  �  !�  �L  !�      H   ,  �d     �d   �  �,   �  �,     �d         H   ,  ��  "h  ��  #0  ��  #0  ��  "h  ��  "h      H   ,  �  $�  �  %�  ��  %�  ��  $�  �  $�      H   ,  ��     ��   �  �L   �  �L     ��         H   ,  ��     ��   �  ��   �  ��     ��         H   ,  ��  #0  ��  #�  ��  #�  ��  #0  ��  #0      H   ,  ��  "h  ��  #0  ��  #0  ��  "h  ��  "h      H   ,  �L   �  �L  !�  �  !�  �   �  �L   �      H   ,  ��  "h  ��  #0  �L  #0  �L  "h  ��  "h      H   ,  ��  $�  ��  %�  ��  %�  ��  $�  ��  $�      H   ,  ��  %�  ��  &P  ��  &P  ��  %�  ��  %�      H   ,  �d  %�  �d  &P  �,  &P  �,  %�  �d  %�      H   ,  �L  #�  �L  $�  �  $�  �  #�  �L  #�      H   ,  ��  $�  ��  %�  �L  %�  �L  $�  ��  $�      H   ,  �L     �L   �  �   �  �     �L         H   ,  �,  #0  �,  #�  ��  #�  ��  #0  �,  #0      H   ,  �L  %�  �L  &P  �  &P  �  %�  �L  %�      H   ,  ��  #�  ��  $�  ��  $�  ��  #�  ��  #�      H   ,  ��  !�  ��  "h  �L  "h  �L  !�  ��  !�      H   ,  �,   �  �,  !�  ��  !�  ��   �  �,   �      H   ,  ��   �  ��  !�  ��  !�  ��   �  ��   �      H   ,  ��  #�  ��  $�  �L  $�  �L  #�  ��  #�      H   ,  ��  %�  ��  &P  ��  &P  ��  %�  ��  %�      H   ,  ��  $�  ��  %�  ��  %�  ��  $�  ��  $�      H   ,  ��  !�  ��  "h  ��  "h  ��  !�  ��  !�      H   ,  �d  "h  �d  #0  �,  #0  �,  "h  �d  "h      H   ,  ��  %�  ��  &P  �L  &P  �L  %�  ��  %�      H   ,  �,  %�  �,  &P  ��  &P  ��  %�  �,  %�      H   ,  ��  %�  ��  &P  ��  &P  ��  %�  ��  %�      H   ,  ��  #�  ��  $�  ��  $�  ��  #�  ��  #�      H   ,  ��  $�  ��  %�  ��  %�  ��  $�  ��  $�      H   ,  �d  $�  �d  %�  �,  %�  �,  $�  �d  $�      H   ,  ��   �  ��  !�  �L  !�  �L   �  ��   �      H   ,  �  %�  �  &P  ��  &P  ��  %�  �  %�      H   ,  �L  $�  �L  %�  �  %�  �  $�  �L  $�      H   ,  �,  $�  �,  %�  ��  %�  ��  $�  �,  $�      H   ,  ��  #0  ��  #�  ��  #�  ��  #0  ��  #0      H   ,  ��  !�  ��  "h  ��  "h  ��  !�  ��  !�      H   ,  �  #�  �  $�  ��  $�  ��  #�  �  #�      H   ,  �d  #�  �d  $�  �,  $�  �,  #�  �d  #�      H   ,  �d  (  �d  �  �,  �  �,  (  �d  (      H   ,  ��  (  ��  �  ��  �  ��  (  ��  (      H   ,  �L  �  �L  �  �  �  �  �  �L  �      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �L  (  �L  �  �  �  �  (  �L  (      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  H  �L  H  �L  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  �  ��  H  ��  H  ��  �  ��  �      H   ,  ��  �  ��  �  �L  �  �L  �  ��  �      H   ,  �,  �  �,  H  ��  H  ��  �  �,  �      H   ,  �d  �  �d  �  �,  �  �,  �  �d  �      H   ,  ��  �  ��  H  ��  H  ��  �  ��  �      H   ,  ��  `  ��  (  ��  (  ��  `  ��  `      H   ,  �L  `  �L  (  �  (  �  `  �L  `      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �,  �  �,  �  ��  �  ��  �  �,  �      H   ,  ��  �  ��  �  �L  �  �L  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �L  �  �L  `  �  `  �  �  �L  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  `  ��  (  �L  (  �L  `  ��  `      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  `  ��  `  ��  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �d  �  �d  H  �,  H  �,  �  �d  �      H   ,  �L  �  �L  �  �  �  �  �  �L  �      H   ,  �L  �  �L  H  �  H  �  �  �L  �      H   ,  �  `  �  (  ��  (  ��  `  �  `      H   ,  �  �  �  `  ��  `  ��  �  �  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �  (  �  �  ��  �  ��  (  �  (      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �d  �  �d  �  �,  �  �,  �  �d  �      H   ,  ��  (  ��  �  �L  �  �L  (  ��  (      H   ,  ��  (  ��  �  ��  �  ��  (  ��  (      H   ,  �  �  �  H  ��  H  ��  �  �  �      H   ,  ��  �  ��  H  ��  H  ��  �  ��  �      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  ��  �  ��  `  ��  `  ��  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �4  �  �4  �  ��  �  ��  �  �4  �      H   ,  ��  (  ��  �  ��  �  ��  (  ��  (      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  ��  �  ��  `  ��  `  ��  �  ��  �      H   ,  ��    ��  �  �T  �  �T    ��        H   ,  �4    �4  �  ��  �  ��    �4        H   ,  �l  (  �l  �  �4  �  �4  (  �l  (      H   ,  �l  �  �l  �  �4  �  �4  �  �l  �      H   ,  �l  �  �l  `  �4  `  �4  �  �l  �      H   ,  �4  �  �4  `  ��  `  ��  �  �4  �      H   ,  �l  �  �l  �  �4  �  �4  �  �l  �      H   ,  �l  `  �l  (  �4  (  �4  `  �l  `      H   ,  �l    �l  �  �4  �  �4    �l        H   ,  ��  `  ��  (  ��  (  ��  `  ��  `      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �4  �  �4  �  ��  �  ��  �  �4  �      H   ,  �4  (  �4  �  ��  �  ��  (  �4  (      H   ,  �l  �  �l  �  �4  �  �4  �  �l  �      H   ,  �4  `  �4  (  ��  (  ��  `  �4  `      H   ,  �T    �T  �  �  �  �    �T        H   ,  ��  �  ��  �  �T  �  �T  �  ��  �      H   ,  �l  x  �l  @  �4  @  �4  x  �l  x      H   ,  ��  �  ��  �  �T  �  �T  �  ��  �      H   ,  �4  �  �4  x  ��  x  ��  �  �4  �      H   ,  �T     �T  �  �  �  �     �T         H   ,  ��  �  ��  X  �T  X  �T  �  ��  �      H   ,  �l  �  �l  x  �4  x  �4  �  �l  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  x  ��  @  �T  @  �T  x  ��  x      H   ,  ��  X  ��     �T     �T  X  ��  X      H   ,  ��  �  ��  x  ��  x  ��  �  ��  �      H   ,  �     �  �  ��  �  ��     �         H   ,  ��     ��  �  �T  �  �T     ��         H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��     ��  �  ��  �  ��     ��         H   ,  �  X  �     ��     ��  X  �  X      H   ,  �  �  �  x  ��  x  ��  �  �  �      H   ,  ��  �  ��  x  �T  x  �T  �  ��  �      H   ,  �T  �  �T  �  �  �  �  �  �T  �      H   ,  ��  �  ��  x  ��  x  ��  �  ��  �      H   ,  ��  x  ��  @  ��  @  ��  x  ��  x      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��  X  ��     ��     ��  X  ��  X      H   ,  ��  �  ��  x  ��  x  ��  �  ��  �      H   ,  ��  �  ��  X  ��  X  ��  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  x  ��  @  �l  @  �l  x  ��  x      H   ,  �  x  �  @  ��  @  ��  x  �  x      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �T  �  �T  X  �  X  �  �  �T  �      H   ,  �T  �  �T  �  �  �  �  �  �T  �      H   ,  �     �  �  ��  �  ��     �         H   ,  ��  x  ��  @  ��  @  ��  x  ��  x      H   ,  �4  x  �4  @  ��  @  ��  x  �4  x      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  �4  �  �4  �  ��  �  ��  �  �4  �      H   ,  �T  X  �T     �     �  X  �T  X      H   ,  ��  x  ��  @  ��  @  ��  x  ��  x      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �T  x  �T  @  �  @  �  x  �T  x      H   ,  �  �  �  X  ��  X  ��  �  �  �      H   ,  ��  X  ��     ��     ��  X  ��  X      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �T  �  �T  x  �  x  �  �  �T  �      H   ,  ��  8  ��     ��     ��  8  ��  8      H   ,  �|  8  �|     �D     �D  8  �|  8      H   ,  ��  p  ��  8  �|  8  �|  p  ��  p      H   ,  ��  �  ��  �  �|  �  �|  �  ��  �      H   ,  �t  8  �t     �<     �<  8  �t  8      H   ,  ��  8  ��     �|     �|  8  ��  8      H   ,  ��  �  ��  P  �|  P  �|  �  ��  �      H   ,  �<  8  �<     �     �  8  �<  8      H   ,  �  8  �     ��     ��  8  �  8      H   ,  ��  8  ��     ��     ��  8  ��  8      H   ,  �\  8  �\     �$     �$  8  �\  8      H   ,  ��    ��  �  �|  �  �|    ��        H   ,  ��  8  ��     ��     ��  8  ��  8      H   ,  ��  �  ��  p  �|  p  �|  �  ��  �      H   ,  ��  P  ��    �|    �|  P  ��  P      H   ,  �$  8  �$     ��     ��  8  �$  8      H   ,  ��  8  ��     �\     �\  8  ��  8      H   ,  �<  �  �<  �  �  �  �  �  �<  �      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��  X  ��     ��     ��  X  ��  X      H   ,  �t  �  �t  �  �<  �  �<  �  �t  �      H   ,  �     �  �  ��  �  ��     �         H   ,  �$  �  �$  �  ��  �  ��  �  �$  �      H   ,  ��     ��  �  �\  �  �\     ��         H   ,  �<     �<  �  �  �  �     �<         H   ,  �<     �<  �  �  �  �     �<         H   ,  �  X  �     ��     ��  X  �  X      H   ,  ��  �  ��  X  ��  X  ��  �  ��  �      H   ,  �t     �t  �  �<  �  �<     �t         H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �  �  �  X  ��  X  ��  �  �  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �<  X  �<     �     �  X  �<  X      H   ,  �\     �\  �  �$  �  �$     �\         H   ,  �t  X  �t     �<     �<  X  �t  X      H   ,  �t     �t  �  �<  �  �<     �t         H   ,  ��  �  ��  X  �\  X  �\  �  ��  �      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��  �  ��  �  �\  �  �\  �  ��  �      H   ,  �<  �  �<  X  �  X  �  �  �<  �      H   ,  �t  �  �t  X  �<  X  �<  �  �t  �      H   ,  �     �  �  ��  �  ��     �         H   ,  �t  �  �t  �  �<  �  �<  �  �t  �      H   ,  �\  �  �\  �  �$  �  �$  �  �\  �      H   ,  �$     �$  �  ��  �  ��     �$         H   ,  �$    �$  �  ��  �  ��    �$        H   ,  �<  p  �<  8  �  8  �  p  �<  p      H   ,  �$  p  �$  8  ��  8  ��  p  �$  p      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  �\  �  �\  p  �$  p  �$  �  �\  �      H   ,  ��    ��  �  �\  �  �\    ��        H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �$  �  �$  p  ��  p  ��  �  �$  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  ��  �  ��  �  �\  �  �\  �  ��  �      H   ,  �\    �\  �  �$  �  �$    �\        H   ,  �  �  �  p  ��  p  ��  �  �  �      H   ,  �t  p  �t  8  �<  8  �<  p  �t  p      H   ,  �$  P  �$    ��    ��  P  �$  P      H   ,  �$  �  �$  �  ��  �  ��  �  �$  �      H   ,  �  p  �  8  ��  8  ��  p  �  p      H   ,  ��  �  ��  p  �\  p  �\  �  ��  �      H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  �<  �  �<  p  �  p  �  �  �<  �      H   ,  �\  �  �\  �  �$  �  �$  �  �\  �      H   ,  ��  p  ��  8  �\  8  �\  p  ��  p      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  �\  p  �\  8  �$  8  �$  p  �\  p      H   ,  �,  �  �,  p  ��  p  ��  �  �,  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �d  �  �d  �  �,  �  �,  �  �d  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �  p  �  8  ��  8  ��  p  �  p      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  �,  �  �,  P  ��  P  ��  �  �,  �      H   ,  �d  P  �d    �,    �,  P  �d  P      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  �,  �  �,  �  ��  �  ��  �  �,  �      H   ,  �|  �  �|  �  �D  �  �D  �  �|  �      H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  �|    �|  �  �D  �  �D    �|        H   ,  �D  P  �D    �    �  P  �D  P      H   ,  ��  �  ��  P  ��  P  ��  �  ��  �      H   ,  �D  �  �D  �  �  �  �  �  �D  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �D  �  �D  P  �  P  �  �  �D  �      H   ,  �d  �  �d  �  �,  �  �,  �  �d  �      H   ,  �d    �d  �  �,  �  �,    �d        H   ,  �D  �  �D  p  �  p  �  �  �D  �      H   ,  �|  p  �|  8  �D  8  �D  p  �|  p      H   ,  �|  �  �|  p  �D  p  �D  �  �|  �      H   ,  �  P  �    ��    ��  P  �  P      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �|  P  �|    �D    �D  P  �|  P      H   ,  �  �  �  P  ��  P  ��  �  �  �      H   ,  ��  �  ��  p  �d  p  �d  �  ��  �      H   ,  ��  �  ��  �  �d  �  �d  �  ��  �      H   ,  �,  �  �,  �  ��  �  ��  �  �,  �      H   ,  �D    �D  �  �  �  �    �D        H   ,  �  �  �  p  ��  p  ��  �  �  �      H   ,  �D  p  �D  8  �  8  �  p  �D  p      H   ,  ��  �  ��  P  �d  P  �d  �  ��  �      H   ,  �d  �  �d  P  �,  P  �,  �  �d  �      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  �,  P  �,    ��    ��  P  �,  P      H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  �,    �,  �  ��  �  ��    �,        H   ,  ��  �  ��  P  ��  P  ��  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �,  p  �,  8  ��  8  ��  p  �,  p      H   ,  ��  �  ��  �  �d  �  �d  �  ��  �      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  �d  �  �d  p  �,  p  �,  �  �d  �      H   ,  �d  p  �d  8  �,  8  �,  p  �d  p      H   ,  �|  �  �|  P  �D  P  �D  �  �|  �      H   ,  �    �  �  ��  �  ��    �        H   ,  ��    ��  �  �d  �  �d    ��        H   ,  ��  P  ��    �d    �d  P  ��  P      H   ,  ��  @  ��    ��    ��  @  ��  @      H   ,  �l  @  �l    �4    �4  @  �l  @      H   ,  �L  @  �L    �    �  @  �L  @      H   ,  �  @  �    ��    ��  @  �  @      H   ,  ��  @  ��    �l    �l  @  ��  @      H   ,  ��  @  ��    �L    �L  @  ��  @      H   ,  �    �  �  ��  �  ��    �        H   ,  ��  �  ��  �  �L  �  �L  �  ��  �      H   ,  ��  �  ��  H  �l  H  �l  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �  �  �  H  ��  H  ��  �  �  �      H   ,  ��    ��  �  �l  �  �l    ��        H   ,  ��  !�  ��  "h  �L  "h  �L  !�  ��  !�      H   ,  ��  "h  ��  #0  �L  #0  �L  "h  ��  "h      H   ,  �L  �  �L  �  �  �  �  �  �L  �      H   ,  �l  �  �l  �  �4  �  �4  �  �l  �      H   ,  �L  (  �L  �  �  �  �  (  �L  (      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  ��  (  ��  �  �L  �  �L  (  ��  (      H   ,  ��  �  ��  �  �l  �  �l  �  ��  �      H   ,  ��  #�  ��  $�  ��  $�  ��  #�  ��  #�      H   ,  ��     ��   �  ��   �  ��     ��         H   ,  �  `  �  (  ��  (  ��  `  �  `      H   ,  ��  #0  ��  #�  ��  #�  ��  #0  ��  #0      H   ,  ��  %�  ��  &P  �L  &P  �L  %�  ��  %�      H   ,  ��  (  ��  �  ��  �  ��  (  ��  (      H   ,  ��  �  ��  `  �l  `  �l  �  ��  �      H   ,  ��     ��   �  �l   �  �l     ��         H   ,  �  H  �     ��     ��  H  �  H      H   ,  ��  `  ��  (  �l  (  �l  `  ��  `      H   ,  ��   �  ��  !�  �L  !�  �L   �  ��   �      H   ,  �     �   �  ��   �  ��     �         H   ,  �L  %�  �L  &P  �  &P  �  %�  �L  %�      H   ,  ��   �  ��  !�  ��  !�  ��   �  ��   �      H   ,  ��  `  ��  (  �L  (  �L  `  ��  `      H   ,  ��     ��   �  ��   �  ��     ��         H   ,  �L  $�  �L  %�  �  %�  �  $�  �L  $�      H   ,  ��  (  ��  �  �l  �  �l  (  ��  (      H   ,  �  #�  �  $�  ��  $�  ��  #�  �  #�      H   ,  ��  �  ��  �  �l  �  �l  �  ��  �      H   ,  ��  H  ��     ��     ��  H  ��  H      H   ,  �L  �  �L  �  �  �  �  �  �L  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  $�  ��  %�  �L  %�  �L  $�  ��  $�      H   ,  ��  `  ��  (  ��  (  ��  `  ��  `      H   ,  ��  #0  ��  #�  ��  #�  ��  #0  ��  #0      H   ,  ��     ��   �  �L   �  �L     ��         H   ,  ��  �  ��  `  �L  `  �L  �  ��  �      H   ,  ��  H  ��     ��     ��  H  ��  H      H   ,  ��  �  ��  �  �l  �  �l  �  ��  �      H   ,  ��   �  ��  !�  ��  !�  ��   �  ��   �      H   ,  ��  "h  ��  #0  ��  #0  ��  "h  ��  "h      H   ,  �L  �  �L  H  �  H  �  �  �L  �      H   ,  �l  �  �l  `  �4  `  �4  �  �l  �      H   ,  �  (  �  �  ��  �  ��  (  �  (      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �L  �  �L  `  �  `  �  �  �L  �      H   ,  �  !�  �  "h  ��  "h  ��  !�  �  !�      H   ,  �  $�  �  %�  ��  %�  ��  $�  �  $�      H   ,  �L  `  �L  (  �  (  �  `  �L  `      H   ,  ��  �  ��  �  �L  �  �L  �  ��  �      H   ,  ��  H  ��     �L     �L  H  ��  H      H   ,  ��  #�  ��  $�  �L  $�  �L  #�  ��  #�      H   ,  ��  �  ��  `  ��  `  ��  �  ��  �      H   ,  �L  #0  �L  #�  �  #�  �  #0  �L  #0      H   ,  �L  �  �L  �  �  �  �  �  �L  �      H   ,  ��  �  ��  H  ��  H  ��  �  ��  �      H   ,  ��  "h  ��  #0  ��  #0  ��  "h  ��  "h      H   ,  ��  %�  ��  &P  ��  &P  ��  %�  ��  %�      H   ,  �l    �l  �  �4  �  �4    �l        H   ,  �L  "h  �L  #0  �  #0  �  "h  �L  "h      H   ,  �  #0  �  #�  ��  #�  ��  #0  �  #0      H   ,  �L  H  �L     �     �  H  �L  H      H   ,  �  "h  �  #0  ��  #0  ��  "h  �  "h      H   ,  ��  H  ��     �l     �l  H  ��  H      H   ,  �L   �  �L  !�  �  !�  �   �  �L   �      H   ,  ��    ��  �  �L  �  �L    ��        H   ,  �L  #�  �L  $�  �  $�  �  #�  �L  #�      H   ,  ��  !�  ��  "h  ��  "h  ��  !�  ��  !�      H   ,  �L     �L   �  �   �  �     �L         H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  �  ��  H  �L  H  �L  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  #0  ��  #�  �L  #�  �L  #0  ��  #0      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  �   �  �  !�  ��  !�  ��   �  �   �      H   ,  �L  !�  �L  "h  �  "h  �  !�  �L  !�      H   ,  ��  (  ��  �  ��  �  ��  (  ��  (      H   ,  ��  �  ��  H  ��  H  ��  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �L    �L  �  �  �  �    �L        H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  !�  ��  "h  ��  "h  ��  !�  ��  !�      H   ,  �  %�  �  &P  ��  &P  ��  %�  �  %�      H   ,  �  �  �  `  ��  `  ��  �  �  �      H   ,  ��  �  ��  �  �L  �  �L  �  ��  �      H   ,  ��  $�  ��  %�  ��  %�  ��  $�  ��  $�      H   ,  �L     �L  �  �  �  �     �L         H   ,  ��     ��  �  �L  �  �L     ��         H   ,  ��     ��  �  ��  �  ��     ��         H   ,  ��  �  ��  �  �l  �  �l  �  ��  �      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  �l  X  �l     �4     �4  X  �l  X      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  �l  x  �l  @  �4  @  �4  x  �l  x      H   ,  �  8  �     ��     ��  8  �  8      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  X  �L  X  �L  �  ��  �      H   ,  ��  X  ��     �l     �l  X  ��  X      H   ,  ��  p  ��  8  �l  8  �l  p  ��  p      H   ,  ��  �  ��  X  �l  X  �l  �  ��  �      H   ,  �  �  �  p  ��  p  ��  �  �  �      H   ,  ��  X  ��     �L     �L  X  ��  X      H   ,  �L  �  �L  �  �  �  �  �  �L  �      H   ,  �  p  �  8  ��  8  ��  p  �  p      H   ,  �  x  �  @  ��  @  ��  x  �  x      H   ,  �L  �  �L  �  �  �  �  �  �L  �      H   ,  �L     �L  �  �  �  �     �L         H   ,  ��  �  ��  P  �L  P  �L  �  ��  �      H   ,  ��  P  ��    ��    ��  P  ��  P      H   ,  ��     ��  �  �l  �  �l     ��         H   ,  �L    �L  �  �  �  �    �L        H   ,  �     �  �  ��  �  ��     �         H   ,  ��  p  ��  8  �L  8  �L  p  ��  p      H   ,  ��  �  ��  p  �L  p  �L  �  ��  �      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  �  �  �  X  ��  X  ��  �  �  �      H   ,  �L  X  �L     �     �  X  �L  X      H   ,  ��  �  ��  X  ��  X  ��  �  ��  �      H   ,  �l  �  �l  x  �4  x  �4  �  �l  �      H   ,  ��  p  ��  8  ��  8  ��  p  ��  p      H   ,  ��  �  ��  �  �L  �  �L  �  ��  �      H   ,  ��  8  ��     ��     ��  8  ��  8      H   ,  ��     ��  �  ��  �  ��     ��         H   ,  �  X  �     ��     ��  X  �  X      H   ,  �     �  �  ��  �  ��     �         H   ,  ��  P  ��    �L    �L  P  ��  P      H   ,  ��  �  ��  x  �L  x  �L  �  ��  �      H   ,  ��  �  ��  �  �L  �  �L  �  ��  �      H   ,  ��  �  ��  x  ��  x  ��  �  ��  �      H   ,  �L  x  �L  @  �  @  �  x  �L  x      H   ,  �L  �  �L  p  �  p  �  �  �L  �      H   ,  �L  �  �L  x  �  x  �  �  �L  �      H   ,  �L  8  �L     �     �  8  �L  8      H   ,  �l  �  �l  X  �4  X  �4  �  �l  �      H   ,  ��     ��  �  �L  �  �L     ��         H   ,  ��  8  ��     �l     �l  8  ��  8      H   ,  �l  �  �l  �  �4  �  �4  �  �l  �      H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��     ��  �  �l  �  �l     ��         H   ,  ��  8  ��     ��     ��  8  ��  8      H   ,  ��    ��  �  �L  �  �L    ��        H   ,  ��  �  ��  �  ��  �  ��  �  ��  �      H   ,  ��  �  ��  �  �l  �  �l  �  ��  �      H   ,  �    �  �  ��  �  ��    �        H   ,  ��  x  ��  @  �l  @  �l  x  ��  x      H   ,  ��    ��  �  ��  �  ��    ��        H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �l     �l  �  �4  �  �4     �l         H   ,  �  �  �  x  ��  x  ��  �  �  �      H   ,  �L  P  �L    �    �  P  �L  P      H   ,  ��  x  ��  @  ��  @  ��  x  ��  x      H   ,  ��  X  ��     ��     ��  X  ��  X      H   ,  �L  �  �L  X  �  X  �  �  �L  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  ��  8  ��     �L     �L  8  ��  8      H   ,  ��  �  ��  p  ��  p  ��  �  ��  �      H   ,  �  �  �  �  ��  �  ��  �  �  �      H   ,  �L  �  �L  �  �  �  �  �  �L  �      H   ,  ��  �  ��  x  �l  x  �l  �  ��  �      H   ,  ��  x  ��  @  �L  @  �L  x  ��  x      H   ,  �L  p  �L  8  �  8  �  p  �L  p      H   ,  ��  �  ��  �  �L  �  �L  �  ��  �      H   ,  ��  �  ��  P  ��  P  ��  �  ��  �      